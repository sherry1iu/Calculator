`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2015"
`protect key_keyowner = "Cadence Design Systems.", key_keyname = "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
T0GRsOgghipdRLEd9FgyHdwknDfUPArww6MW9m7Mqo6md6EHAd8FeY7rvzjgflJoaK7VDbka8w3l
JJYBsfvGhQ==

`protect key_keyowner = "Synopsys", key_keyname = "SNPS-VCS-RSA-2", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
XrzcquAd4rHB2VHaZRwHuQPZfV+8wq3+lZxbyHD1LCFC99QPovZJYMtDYa/yg1gPkxapn4aEwvnJ
JdrZIj78vYbneHK8iOdU6YUq32eoEPj9qJadpln9ArXgvwHQOW29IGUnus+SYnzJm4C69MgMEhXL
xrwkGL+AF5md0PW/1FU=

`protect key_keyowner = "Aldec", key_keyname = "ALDEC15_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
sSsUpc5lDn2J56zOv/OVYnZf9WGYxQs+Cm6DnOsVQWnCjOyYAnhOJUAovTE0YX9qEs78fecUe2sJ
RBIEaZDJUyNz3SN9TgDRduNi4ELDhKDZIQ8OXKX+MpeLMgb7NKLVBq9dKKZnNGxFqS9UzlQ1ZbPJ
wtYnztVwsr5JLqifp/St3X6cqlI/tOKzEz8BUBInVj01760dHe6E0KRWhTfzVwA0r5luCErt6KcI
L5+jxFwyjIF58WSjz7vxXdb1r9Whs7McvEjKJBwWvEWaAJm+ufb+OGca96Gp4JHKbeEWgtZqBPc5
52bYqqckIl/+882LND5DfwAsnuxeAr3bOpcbfQ==

`protect key_keyowner = "ATRENTA", key_keyname = "ATR-SG-2015-RSA-3", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
f2nSztJyGK9Q6mZ5UFuQdKIPyA0ZEtaEqJLnDF41ssm6WJEsAImz+WUhWNvhib6CO+paRpQ7jlkO
vPrdRurWd5hQMnAXjkmMWJa9iSbJLrC+GBBBq8FomwBK3/88d6MMGVz0SP8lO1C+J1+G+sUqqbjR
SkTl0H40s2lOCwJ7hjvFL6M79TZJX8Uw3IM9vAdMTEYiHGvMLfo+jO7jG8NGObilbEh12fw4pNYx
yJslmP8/maC1eh8FwBX5LkC4eu7D+hSR/vjBj2ExQ7oOO+o8wjDWzFGiKGVVYUsRc/S0+LMbg8l8
WjCv2Z8jTVWHnin2uSHhXNXVyzXLbJPy8orklw==

`protect key_keyowner = "Xilinx", key_keyname = "xilinxt_2017_05", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
QWcidyxQUP6jobyvbo9q5AllRhQQP5Htpzt6K17DVIHA3trJxURDhWNbK/uW/5xkyNMCvaChM4ZA
y56MW4Q75zv6rV9nzlGd3DGQ4jneunDQTixU2/Y68HuHOQ/01lC9gupEHJHTb3x+nswmMOa1mYw/
hYeaGs0nh/yuAx2MzuLIduBJj8IiwHScUBzDxriHtBHFoiJ5qSdPc9gVPq2BTxlv0/3Oa6TT0RtA
wjVNjAiu5DbWsSMy8A3pB25+ALZFkY2NYitVvGMqr7AElYiejfNU4mRyqBinhmrm0cKJ5rK6Cdx6
Xvx41Vqu8+pjEMJmkun6+qgwwyBy11VPGGC67Q==

`protect key_keyowner = "Mentor Graphics Corporation", key_keyname = "MGC-VELOCE-RSA", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
fQbPowMh8eLH4vBHBAR3g47FqoGtEZXeVk32KA1WcUzVPlxfeqTbgGgUY0N/AVptX/s1fjEE1fXB
5CqnZTRFKSGaCYvJ93kkeYnhlDHSjeq+PQrzjd1g5OFfM3tR9IPBTPV41H7dEPO97UFty/xNo+UG
jgnul8ZHraLYJ/G+rPA=

`protect key_keyowner = "Mentor Graphics Corporation", key_keyname = "MGC-VERIF-SIM-RSA-2", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
lBHIWl/b7qiZD6hFKjExtOXdaN4ZZJk4FBTVR+jv0cSBviEC/vUr1AQHzNB/b2XH+UzYrtQK2QkD
Li2Nq1jjlkj25Ir3Vy8Mh+DNUDarvOF4o2bAm5P96O9jX/WFFdTvx89qdIrXBNEbnqroPaB0bHUS
f8zIAcScmoqB8t7hezWm/EOngHLlnOI0klm3sGxCdg+q82FnBXhlDpsTW/sa+Xb64oqKWhhrM5W8
1jRVaV7ERFAHXhHDUV6S8TjoJfMn2BMp0sHmWaC+TftWvP5wp5N1k+dYZSsSLT+dcPAZfLwiG3b7
QqL+r+zuT8tqI2U9unVKxFjDnKUpkpg+xjhpgw==

`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64128)
`protect data_block
9nFsk/ryzPn4rw4iPal0Xm545rUYrN5OWYT8eiXch41NWdbzaNq0tS92PcbGf1jBpOSeabqOWa/J
IghU6FbpDW7a7DZrxxdo/0HnpoXhcskvj1OkJ5QG+5PFRAyhXp6+QvTu05Gb3Fs9nNMHLo4J4wkS
Gekz5Lggfk2SVM+X1wq3jX6lqQmeIEbkIrpaChI23rMjRA5I2Ld6LexeYa5fzgtKXTryCwHfyWgl
BzGXrKtCsg/mqAzjP+JSRIA7STG5EpCU12WJxGc4tNUzectSocyV9CmtsXXZ/1P7NgPo7tpVoT7R
HHlxyVJTYSbVwMb7GmEVkgDoizNSqERCtbNYVHbY39ll0ClUNk+3DteOVP0/sh1/qMnHzl9CTyVl
jG2PSwoMRVO1djFh/UFgDyYcsLeszFLePlMvNYQxm+qf7eXlYc84XRT/0ZRS8LuzkQuXvN9ZVQaq
Q4RfEFU+1iF9ift73O3Sm9JXg4iwoeInNy70mP+Wyy3oQ+nuL9LPZJeuvgTyquBSzejzL+YhVSvT
ydqXkQLJNaXRCkxVSekIEmLSxgYdR8n8kAJygn0NDzTcANDPZVAb4alk/upSXF/V9n2s91yiw8hl
sLBoCLWzwhmSuS6e3NF7J6kWuQIoRA8oNRwWDqK+o5Li0V3YFjnxjlNU03824r8pPURCcn3yFz3P
QpU+B2NWDa1468pAJNRouiFD1l6jJ4XjZdXkWNhExbpsFebGr873ygHJVJSyl3wNPp3YsFKoLOK+
FMuG08wH/hd0Q1kwJNTfz8wXHTbeUDZ9NMIGHV66ZTrwrhFlvl7l6O59BtruQ1DnJFf78ZzfOebc
271vIlTua1PF7cgsDbOv88LxwOfliFFOQr4wkOfzvaI3A4b4p7N771+Nasbt/jqJBYOozhVRm/Py
jX52DBmMIR/KH7thpe24d32Ej0333OnTMmq6nNMgjNq8SGvchJWOmZZLQDNleMrXzjNoaxrIIuMt
lRruDXty4zFUDfxQapwjio7wEXqaVeiWZy3+bM8fbxz2pF1uGMZRbIfYpOPQkkfXqO+5T2WoZrTo
ki9KShPSKTAKSXTJt2pjLWx1YB676Nsi0H1KJgfrarxNev/Su1b6S+89ezGu9525nHBxgX0iyWHX
OU09uA+h+gwDdGyNC/J8dIYtYebT31jX4r62TiotJ1PWqLuv90s1uhVr85MO1FyiyqzEkZvHF+BX
23ldBbm263yz/H7QrfhfW0oLVdV9FGpWQyATCCcvoF6OoGJB94132VB4PBZMS6Y2hdlwTuYcZT+o
cjYqmszhgQsRelVT3aeIqIPc5MGw0HL5yukG+OteX1WPOXEfuB+uuq4qPnV1pFQjMPQU+g/VQiBb
4tJpaI7P1HZj9KNqLaudBdTAx7+p5CDxiTACu5RwPWKDgdDVwdd9hUg1ZPg9n/TqTu7IMWBoH2Iv
xtUeaegzETd2LfsrO8n4RLk26bWZAQM5mj+uucFBd4XzsyCzUwiwbz9RSLouTYaqXb27Vq+Syc59
sH7A5agkEGPyR3C8ZC34LlhiWVkEri1ELsPnbDQmYkPhZwRowkkZ3gsHYreTjA0JmMb9HVLQmqxl
o3LfVq4mGJLa3PEXY1IhGHo0/P5LmiqxUrMJK4KawZk4TSqZHDqWNk8WN+xlfLoPIOHmo9bMquP3
ZqNFgk9jLu+olCnzqtDYyy9LJNWDKco/qaS/I83Y+lMc+TjsmtUeD6+lCgezwGSLnmsJLT81bfcr
/sqRBGSk4cKq9UKprXaSPEceUJ/vTGCRKXPmz0uVKPXxbN8HvzhlK5OwgNwALB5Z3/k+DAzam3ry
6eWFz88uGtZta0tFJcPC7PEEZ8hI87ZPj2sUeDfpQvp3BPmty/TgW3J+vsV6aV8As9TI/fxoQ6Lf
AQgNyRjXxvSltCFmqGnjlN1QkWm3rjYhzetHrXnuqeUCuHOwsGOJ4VCWJtW5bW39Dg5HS7VVgRp6
V3kxM9mjsWwnu/2hEggf9vJQAEoE/FMzwgqIY6QDXO1c58Og0AUZzDWMe8kc9D/nHAOZEZAGUL8l
y4uqVsLQqhZ1aA6VIY6yshf6Dbgiwgg5ZA9HF416qazhKlaJ4E0HqsJnK5TelmWZz3QYmGjItvg9
8AcEEKvnG3b0qMU7sozWa8SZuMqfcdJ1Y+InqlNR0H3liQ0mzlozkmcc4Eb1RS3hA13/LmA42G7a
DgnYKlFg3mxyvUEdoIfAK/hsQPf0s0s4oTDmxpXAMVmfKrRjPMnyJ7o6hzTv7JYnk1BHYscnEPgM
KOza8cQ+8rHNkEAgnTnswVHZLfobB6HR3f2oNG4ILak4G2uYnhW60da3nyLWLhnkgY7VogxT5QsE
ogTuiMt5k3K9+gti2Dh/a2Pp/vBkwzUOyx5LDo5N1JDR6AjwLNRENGICJ//G/Affmpf+3NddkLPP
wr/a7oBTsKMn2kzMi15l5wqcRwCRB1DG1JHAWK0956CfM7s8E9UVthok87LpsQnW9fjDckqwF1Id
Vb9hgQOgdv3ygL4MCSjUPQ5wV9xnzr/CjUrzCjawTTtn33VvQmpK3Ir2EwReBgE6BExZbinZNm46
i2NP2BBA5QKmNwSP3QeYXR7JjWmmylYJ4briBt/ao6CRtY8pijkI2vd6KJe2+2RVFs5fMw9R8ebS
hDTCLC2cJWx3eez0QIIVLis5f9/KQGWj0N0EQyKFCuuCpCsU6pHNhIhAu1RPCLJ8iU6ufzLtkCbk
jPTDsFNH0TTeFdAktf2ZdTpcbIBVTROdUd2rtBTzL2Jv8kvnIU4xjVy/hhIG9TyyYj/M+bgBvaE6
/kp2/864fTMLlNl6SNckAwiA6j1xa4GDdtMOPQ/vWNmuZlOA/6djC9FpBID6wExU0Uk33DVyH2G9
fBqm4ERPwdzIzPhyy/JP770HEYPhqab57liUECgBMBM0193+esHDQQwYywcwHwjk+G5WPQUEOQSY
jRty8o23VOZHmCr6jHm2nsuE0T07dakNjJv6mRY9HONqxRgpztNcV7NXizsLcfYkUP9do1D7Kh9Y
Gwb4B5Flfu0YRf/G9NAJrPmTj1+YGin4KOYkW4b0zoSL7wJqERSuNZm8FJ5uMNzu6YLwmfsJAXog
fe0EOXuQkSUms9xo2QAxzzEMFmhH6k8WZXQNvtKskPnjLcF50C17c2cyRke6g9xUhzw92C2GyZH6
M1ALmeag5XzMRDoBk9enIognJqHfhAsLJSTXPaar4se7QDdWrvd64G4HjilN+5PwTV0GmaBzV0qg
SpA5MaaTY8LbHWl5Qd3DSlgn+6uStW+jUdNT9mn74atIIqfBp3KqvdaE1Iuo66Rn1JQM9mUsHz3o
BjTJm27ZCgul6fbmFyguLwBOW9qyM7Uk0eihZ3DchEM/1h+rKYZF+MNeNU+MeQ6F2m7D0ii4iZgG
pMcPdjekuLkG7IGOt671dps3KZdXVfXnjA/qll2e9ohvXwOlYTiSOAqwf9bnMZm+lYMXZf+fb42S
pvf+0UD94B8IFXmkzNa6Cz8MssKbAfm2zEJwFgGBXv1IZ7hw1aJM11c3lgYw2Tl1I1O/SRDjHPCN
sD4gkpHVhfQ0zbtHBEELPUGfEMWFseTC6RRbVB62D2B+lGP6I3eGwxlkbY+OrVGLfdAsgwOXDo7p
7rmxBUdSY8iFg2ayas4IBAAV9f48b31my2qLBdP+/k2j6c+gCp5PnUTUk9EtLKUNayA5tyGN+tbl
JeQ9fEdEt80s0UvOsTE0L11NKgkc2ZrMF3eKdJmi+JLui5zktK+xUkk+KF3rerHJnjM9kQDj3fkb
5aPntZ2EtZNNr6mREDTU+fINA85XdLdtZ3LOlCK3FYimxy6CxLZJT7cn+1eQcm2VwjLmhVQCUAga
zWPPxc7Ikl6Gri87SZiFd9bmCjiDCYIpBSF2IYq7t6ppuxLZLmArsbf7rLfWzjOr7NgWE8I18vfH
98F/B+DXs9l6h60SgnPo/V62pyHyjsNxzM1tIp0rG04cbTJ2oLlcPvj1ed6HEafzBvrvkDQ/czog
Hi/OwkmGWTfNvTJSn/C8bnH486+FjBP5PTnxA+REyB7zv/mcBva7Q1KHUMOm/VvWBUCp6dIvKMUB
b1U2bonhJSCqQYInRFigz06dqAPLe41pQZ2qBcGNtzXx/ncuHaWyD/dExKLtSbX5k241ioujMgWn
N2AHueTqBbt6jZH/8sr2TvyEm55mBXzTdOhD+Q1QOv/B9ifNmVzD8KbXBiJKErp3CltK2SMSnukk
Mr9G89mwIZYI3nM9LC45ZqdTB25HajkA4WPJJVF6n6/m90mrMi4Wmx3/qo3pqt/hvnfpUeMI9PjK
29+XU3AIiMY1w2ntThU93mzVG3OeBfvc8LkYqOJp8jNj5/kZDqmENRH3wquTkcDmlqlRtMax3jim
CtRJnfxboI84ejTk0cxfBn+jwhTNg/yf221PTiKKttgL/8AW5l7Obh2gw+oVFThhZ/4iKW3bMT5b
Bez6biZsozq5D6PFYgI4hTv96keaPB7//a6a/T4Ua1iQu3o3OPgc8z2kQ2DqvHMzUxUtnHEdW8kz
M0JhaOKxvdAE9OGnEVVZ9IHihyIz9m0ffGENdtIBdVSCzkekiqraV7oQxh4WY0g/5Ja6Qr7PB8wF
R4VgCi3Y6mzmZozk4agKAFRRAR2y7fQAHXM4PtKEVpbuKmMnBR9katvtUgXe0Tw7Hg0HLGMGTVcS
A0EJERL3B22CIDKuLEqvWdtri/oDVHN/TB4l8hbVtsJhPkeuBsg/7g9ZZ3jPmXrm4oeIAX+OvgS0
EEhh1ExKpqMWp9R0C/SoCyE5aLIfo8jvE64lW3R9V/wC7cK4CZJLVaWWLZB0jTe+KC6KsqlFp51Z
MVIIYCQ44sLZP3Y2TNMkIYMw9O1klm6Qq9WA9axJx+Q8JphBAH2QmaTI33pAYl83efP+9nfDBzod
0eHBPZEMslHBLTJ6qPVgvAmUYgkH949QZPNrrmW7MUI+AXCT3DJpg4ZBoA44gUp5XhostsJaUxke
fhkYEXTVV+ft7hWOG4FUFiEjwnlfFhuDtNvP7ybMemof79Zmi3wqAmbBQk7z2M8rSYLO5DHrZYOu
Nud93vR7ltXvSeWe2bPEF67xAfmBheLuSCTqTpL9H44sbs7TW5snj+WohK+A5Z/ifCWmQUjOZX/L
bGDWrze+iMgo4zULg4Ebl/xb4jfmXsfu+IWBCX39Ew6G/OfW65LWiKv8ZZ8LMxV0eIeP9GuufqiK
s7dNwAq3y5ZPyeUDaq7dzzfua+daQOQKHj5XYypJ4JB94nKknL7DJwvGFyARDK8zR8mjTrbFvOP+
ES+XT2aFbOivxnp7ueBUJwj8HypPO13TJous82nBuOJfnQ9H6OyQ0gGkPnmzQmZctPkwdJlEYiWv
kQ5XV7DEEvIAZ0aRf7fPWNTxo20cyZNEsM998NnDmW9Qo0EPMxazpw+9d2grZJiup4vmoxBOA5lz
mpnBcBJAZISyyNvPFvqxYza8zG1ZGp3Fm08tA4iMLiVC2pHI9dPxgYaltf4Fw4NBs511xJ8lCMUo
SsvaN0nrPkO1y9kgq3C7XLzDoH+we1aS2XoN56W5QCt7sfMpxpBkoR0BRYXOWHf5kgqJt72EsgK2
bSwHoxbxPR/ZAvLNtCrEbozzkigv8znNlCiHvRJvno6OJjUnPJlCJI4ak9beqm9vtXrIH0B3unfs
IgBYgulUXxDzqVQxqvHxjEVhA0EYN856wZBgziveJGd8rlzem18QTLsybJ2aw4a+aZ1mU5/qeGMR
ZO9QDZCl5XfvFSnbw8zrW0MsSKOW/uE9vS4nbIxVC9LGNBQcne3/7ySVe3ocdW0tHKzNkdSc4iKE
2H8tA/LX1vxFogjD35sLHPMeFCz8LDKkN1H/ZTT9+0cQWTXN1ZrtIXivk2APXj8esVQJWEKNGTbG
1B3/kG9/sy4uPEUgCPDJFl9F+/Qbss6qe0cS0IF5Zyf4JxPdFEtYxeBU0pjgxS39eFWXBLEGzxVO
rebePfvy4UsK6aHWLV626h1bY9tpjfZO8gMp/UAYaUIdk+CD7v+JFbrpY7tFGFJk/nybd/KlsoCK
nVEzl3fuJwWe6hxptDLiSNyXQJEWyTk79QRI67TLedEtKCzQSJvLHnn3AuhzMXame2glum5bW3U0
ZOhfTBdkhyai0QbYP+lR6eAkdzoIo/kbzwy4yKG2ql1AB9zZF98gMa8Pq/1C+4cwQ6RNwLQRbwYE
MbZqW9LL94xtAq+Ff5MKy1IVrnV89Q58/4PyeDj8IhzgVudaFPp9ntvErNjVdSLCD1mxxXvwq/5y
4+n3Ym/UWTkd8BYChE20xMcoXssyoF4jf7XEe4KqnMBLaCU5A8WgmasY9nuX8v7PUN8vbEjWYps6
BCTZs/ZTWymO7E+48BGF+55NZcMXXyeNS+z7hAX6w5Ac1Vk7ce9+NrU4ldP0lCLicsQXoCsnZD5+
lZnwKyuz8m4eTZlFlz/exih4Nbw3cC1t+7KiRAgn46yDQolFbuJ0OAwSh2oX1qaHdmybr35JCXZ1
wODjZHP9L2FA5orbjqRB1RMsywDLnasjguhUo9ljvaX6WLrM8Fd/0ojhaXtUT+a4nMV4APu0eT8K
c4LRl+5lUfMWAXWFETB+Ehy2HtSWPMetfDxPsuaTyoo7Kldh54rE/PdplGYgvwCpYVSBTUNIZ8dL
Ktc/uoW08omFGuWoaYrZ2zkcJZ/bFY0TfmBqghBJcLR6ApjRWUCpEQFmnyZb5xpMeuUMB0k/oU0l
O7HzTj2BMqLgZDbRWdqBMGTelsVLr0HuP8IFpgV4yLKE/xZmENWVFmiul4cIEiI5mMfVRrAGLyb7
oQMPRKzRuF7qfufiqJg7oQ30WownAT6CN394yd4Pd9ux50DgEAalAfMO9Kq6lRcei4sYhhFADGsN
OR3qQ24ZfP6b07R0soxNshy2iNvHqMFuRrSpnm7eLSOvzE5EBXnCng9nKsiiGv3PTar2FOGozexu
w+NsIwEol8KAN5RSDkFfQtdW7lS7RmK7hmOQgEa+WZlWz+AOnhNd7W/vtTbUtifQQXWvUzH3AX3O
YRI798Q34fHuv1d/Fdx233vk3eDPlxhv4h5+1o+6IEOtWtiVVmilnwsbuSUM8AVacVwpgRFCDBLv
ZaZmBJ1eWd/1NyUeHBVLiaGWTllizNLhTL7LPd4LoWIyFFZkXOSFfc1PZRcDm9novIyLSD9gEcn6
a2NJZz3DDgstISSmj/hHEu/LfBEmNCln6ogqQIXzkRjmhfCrZHZH2OlLi3WJJEjC2ezyt2idXYdW
Cms51tsjC9CPdjLXXoH5kp+puzW2gzXcNqbbdHG/jiWKyB60RnwLAYe51pO1VTCjAMm2IfT8y9h2
z/vXHXWJIRH/BINlf/NP3Gbsbq/h+OTi2WpAoTP+yKXGUBA0Dav7aFBzHBzxdNd+d5CTR6It4nqT
dkHRP1UUYHAgLnnQuMob06xnp6bgdUlpMzAfH6hk6YHWjcTGcWpHeLVQfiyrbs6gJOZIavLIygmJ
qKnqIzrurmM49cheA4zIaZSwJ50tYcChEEL0dHNqTf8gBT4XmMxt4ORE7dBBsvFQ9ZmlF3W/ixhz
o3HX7nNfGYkss7L5Op61QWliXPWK+DX4mnmPptazWhxuHMKnQFV95F2c0BcG4g6ydBesrNK+k6Wn
ui1B412c3FmTgJVgvuvG0OvHIS2wssziHZWMF0N8lSp3a2Z6U1W9Z18JKwgOKwU9y60pHLSc+esY
X8URS7EClCqNDL7v3kpDSvw5QYiIY9mxrZjSolEiStZCzToOoRrWWFc4U1JTu7t9XChuXT+poWAg
/r/UsFkbzvn3+S2M4DIpIkhKF6IWZNafcyOzO1paJFxtH6nDc9u3WjViHM91UNjy7NgTvlbBXaDJ
HGxdks8MIfOjZpWW4lEGjpwj2alzlYNvZh47/IVITllBDTZ3EU6D6trQrbQLhD7ZqU/k2Phd/jJZ
fkswCZWum+G53Le7+lD75j03CuazUuFZyBpGy3TiHX53MnRdH1FV7kmGfYQQhNGIk9NMhCSEm7ND
8n1EwI1jyHLdCBcSwkbqm25oIZv1mML0nGZakLjt4i6cwa7Hpdo4jbuPRg5pLYYJEBZeBTLTPpfX
I9VBZaysu6Q4zba0ABtWZWkmMbpByn+3FQwQ09KXeqDqz1AjjJkHDo3Rvx1q9Wjj1C74m6lCs8H7
mS//JYRe8rUfHWdLuDwcIbi5QDnJ9nwrei41Xkvd/TnsKKrn+yCLBEtwP56DDfAczE5JtuBeYuwB
YaP8N7vvbGCHXHZA25IVkDWpvPOBk2k+RUG2k+g1yJ/iQ7KUaikOaUXV+tgFebaAsouCFpQ8O2cn
mGBwaRyk1B6bzjYGzWsqoB5VXWYUQZ9qlFC6mBFg5Ox8PEq+/mJgYoNosHC8zPpAiGZO3a0UwaMp
gt5N3C0guuLctXBEe4TZ/Fyw4OuNQcBmFx2uTd9UeYbs0rUffBaNvLLBIY5bIOr5+cHeG5nfdZMn
vRdNU4Q5pJUtWjCiOWQ+xXs1ZYEGXJqFDRgKjr2yzqjvEK2bLcegCFjvIu7LnUkBsbyujy+GfVi5
N6ShOCv1oec6RaEhRNY6GhDE9F+pv4pVMNtD5uiBRNheFfoR8fDudBfrSvSJfPESwqRkEyviUqwl
QNDNpVuTU6mK2VpKQzqzfANRQTxnvDFFiIM4YaEkYvCO1ItnEpXk8stxN4F+AHyn3IXVQvTvRY5H
K7fX8wKswfnSwvBOBf4Q7hNSUY6h0lteJYy4MoGICRabGRhb4pf/8KobFPnQeGNycqFnWQQ84ZPV
UmIM3iMW9UjD7s2Z5ddZPkqUlVnxSsWXl66WHH51nlJZOHwtrZM6krXn4Yo9d2PD/xJPQYeRZ5ZS
Qf3mpTV6Zb/uT6Th7zRvdQ3Ib4SCWPMrZMXzByzscg+0EdGgi+1Lyo3q4vgJ0VNKiL7tMCgWgjBi
uqw2w3uVu/aHo6L/KFJ6N+pkBkT0lCjMtnQETrZD+mQ6CQOnDTgu0JpFtxMXaEWs4Gvt1iYdKi9r
CRlXYxGD9vcMZOY00VRT1ZEyK1zDGVWpMnolcFGs0kPpum3rNn+KVvwOKk08orDNdqqCTAKgSD/q
K9YH1dPozlNLSuNcVjgJwtb5KtYZKaf+SCeApOIbwz97y9fuF5LTwfzZs7aTgKzzlsiYOzu4d5vm
4kq+d0+CQnUJgwT1mNaX1x0G2VWlY6Hl4929Ehe8S+wGW2p9cBtswgW8NSqGOllCRMQik4sIKM6/
ZKmIDqx55cDnVbNladSuZr7vcYsCifyVC29xDxctEhRxKbaVPLXk10XZ5mrDCR6zgqne3qWJdpmk
xQw0wrOwCvEGdvbtyZv4J/jTmgGVtoxmjfn+Lmc0jiwzgbAlhqiNYiO+5S3e9tIgFQVmZXK/Q1XP
HIqJy20KQZOFW4VZ1TZ2yR0lgd4XPJjqaAalnbGApZ8jpuhIklNdvx9qOSqd45gD8LUZgj/nTXJB
QRUjLVuBXysPULVxVDZF4+fF1HNzBwg4XC4v5/N8liyLBepOfLr7Yc1XRSJRcDWWPUY1JDr8iSMR
znz1/h0pvgF9VB5qNmSpQtYzOkkQ23XGKf5SZ5EZGiUv26DmAUY77qud3Li/DRMTdCD8SRiKtc+c
kZi3geTB4rPQZTj08UcEUKerc68HiZHEVYbiLXGkuI6OeXX3TRF5uUzR+F3UmMulm5HcGHUfbF9J
ICF7gRKmfu1Kjbj+dK8BX/kbHrrqfx3UL+SPhaNsNwUGv6T/gpQlq1Edu1G2P3brtHtqagaWSkIn
eMraNLTruVnADrSyNfaBQMLI/3BE/4Vu9A1lY/A3UEhhx4ptnEyIg/br8s1bOWDcVTJo4ML2XbBb
Q6f8ntDWD2qHCZOf49CLPXYXisgubeBCChj4virINH536G69Nbc/1HcHCngZpt3lvXmByaPbllSY
kK9Kg5/ZUtHKg1s0jZYPLxz1wPmi9nthkcK79veBvqonBgl9ap4HgjeZ3T5uN8U3wgA982EG8Kzv
5zlHnkCGq6/jY7WkAuR+TsoVLvbP/bzG8IilWh9MyFxdSw+3R4FNG5TZTCltrjmCu4yF9Cm8u8RK
vlK8ldvqM2Zvi3NQ/YI4szCfrux8sLFnMllWU5GMVRegIOmLUQAk4wA2c+i6n2hWhnQOsdb8E3CU
j0XTNtOq5FoC008kge3HWuln++vWTqBWkRc9meT9BZxKDXV6wWZM+HqpEprcG040TCliqCS/WVD7
A1BADbOive57n6x8PFtk73l9W1hO+iB4uWfPQx7GbyISXVUC/OjB05skwgk22BfAaysxTuGkGuwx
byeKN/FRVg8cG8USBTHE6pEn/SXVi2PE+EIJM40UvzKRmEbXiTDAkTMnk3IV8TWwCAvwq5r9yJwd
kA9V3vVYxUK3+WtPp/oYa7fz/YI2XEQ527S0Z33yddNMRyxComZC7sIf0f8nf++Lq5LpnolKFm/j
p4OqP4n6i3/MuwCqbgMgplmNOJUOSCBjHGgc/GKDew2SN7r0LiP6m9ziLQh1x+PV5DdNFhH2FRGn
t++nL6Yy8eqJUFlNft0ZWM+rMQAPCERnad18EN/yvJBaZP8/Jds0H+Dd7cGDX72Q09OlZjJZbUNn
7sRLjQgjqV6n9ta6F5EI5tQfBnseF1hupyE0eB3wrmMG6S/nkivSxcrmeZKR0mUUsGnWB+NtW30/
/loLVIHubRWdsmGFpnkmU31eGqtuZmVz3EnSjzBl2C/45u6u1AYtrDL3R2QAOnE67Q5qywTN0c+l
9jUTS2EzmbAeOEH5cil13tl5eIMw8osSMFgQ1x+tq67h0qau7X4YopXjivzpHRWCUkEIevlgwsp/
UNFhQhRG0YYLtR4xJKs8jEKsyE2w0Yp2OKNwnq/qm//yupcN7CNrTXkpqYvJWJIh12mKwKgX9Xw7
B5IxCZXwbm/si/lGyx5C4lxS+t2+kfd9Yr4gd1JH9e4G7QPDvjtkc6auWosxk8BFFkNFqC6wko/9
rMHyheh4004jsYvBehgZ2/pjejRzw4AUWyXlwFXd2F/DazPu+RjShQMXi3I04A57aQE5U8fWbKu2
Q3mp4OF8GntpvG1h0g9JFC8uq6OmA6MciJkimbrn3Qjhf/kGrwciJKFOsh3AiO3Wf7MVkAWinF4t
94CHVrnO/1kM358aWyjt7o1rLLhY8o02sh6f2TmQZ+RzgMppmTDuql8/7Jgy/bv6SKPQ5ig1hAt/
yQCYU8e994yWOruu2SARba55oKy68hkqoLRPRL53HiJr4NGFQY2rJfCIbZ/Ni6dvObUWX90jdzxd
T6L7NmeLHX3poA/mel3pY1Y2LnJzLC9n+yBN+guOLWcaDuK+moPWNmv9CbOH6VUodUzJeR+I4HZF
7z60E4rgJjBLkerGnzJMMnBHDUP+v1rRiJ1D6AacbxLox4DXjdjq+X4YxwN/IoM9wCYnjJz6dFhc
AYEZdpUb9fZIvSvYGRTgZlhaKbyR5+Wwtwe1hlrTvf6efzMxLcI4qgeGzwol2mox0RxiEm8lsRAw
3KJjV5+EYDP3s76NW5R2fmHW4VQL0dyr1WvJdUON/ZfpD9ei07aJDaPuuK9HPRqk27+tTeL/AzzO
RizT5DhSA/PxJaKF25igqvk9meZBd7EzNtM622u8SIHnxAmu2g/aKYpLK7erXrDL3ijjkmvI9jJs
Gw9TCOVl2IWL1KuL0uzQNhGQ0FZ7qJ6KZpPOJD0ftBk0uwDXs+KMAvF5GqSPKDp55WEW4GwRMAw0
NAamnRbT01TWSjSz6RjwaD/AFq46p8IwEW0HIkpw/b9/FUIg4SBRJFwuNHVs8HqulbK/necWa8rO
QjCu/hnu6dGt/jwZroB9kmA0u9+VGzk/IB6PPLojWZOE/yCH4g3KzIWGVSv16rgOfuEKq0fcdV6N
zgg6opFkXQjysJ7FVnR37ROWjSKMj6PHJbNvcLJIXIF1hjCth+eH8hcvTeosu7q2ynJTKi/wIdU0
6pJE3AXHk/zIa0W9EmqWBp1+p2NWufd0BRsSoueulNxLTBB/9ncTFK92Ctfg+bKZ6XIR74tIgFMt
lS5qsvMIKk2w5atQ5GPu1L8xeZ6eICxR7H0o6RzLuwgqfFGvVyWPHnL2tKheT+FfijiO/sFbE2DM
+oN1Qz7DA/3P2Lm6Wdf6M9eHBYR3iAua8zfZLPUbfUm8Qjtn3HlYceuupv+skKoL2b5otOhS+FVe
X2s6rIGKeqIbF6B7a8xj26BKXg8AXVG1UqxXMHLp4uYb0l54Abgz4PWlTNd7/wKkNV8RmDW7+y7D
NwuFGIMKZodbe1gltaNgmSBH4PWiJeqM/xMT0zbW3suD2ytLZ4mAPJj/f83sixRobM1zgLcm8/d5
lJjafJ12EsbBPnqF07K73wvm0y2Q51ngY3scpzZiF4e9y4Sz9A+d4jIgKqPF5gC990B7Q2xOZ/sI
bEk7q3KmrXok8vC0X4OL/IbQZ/X5BavyR29359Obm5JWZNHK7ApUf0rkAt3iZMGUKvV+3GV0/153
Ps08JUKZ55WR7ItQs/tsYAXbYIKYXXkrNnkJmw0uPvhZMcixUzAc0QJq6ehNxkpYP46zpsKKFtY1
CXmiL5K+oX2wKSVuh9uRZh8YlpdETTdqlbFi45n35PznWXkY0P9CTcoxj2agqTd/Emzm8etGakkw
midYaKLoyd/uHJqVAoND0uIaxS9A/+CcbBZNUCqxToHlHVs0ZYbRGM/3oMDAf8TX4sskZYiXEKWr
KQdhYz13F4rytYlzlWsD+ge8lV9HgAc7GmK+1B+sYVmzeXIxrI7pBv1u6VgKVb3rxLJcGVHv8rhd
WPQacjJ13F1LU/fnp5f1jgOXzMxrwx5uwZgEhCzqQwhH6Dsu+D9fLpRxqmMvbunq51+snO1Ssjg4
JZLPKLfX66/czdb4H2U7meEcUG22MgiwtRARZVaDvVnPVq89LNPXnvC3xAwhUQaQCbyRlyJyFst2
k+kn+T9abHQATQqKCloSdP0W0/uOFN9WeCVTfskfFJuBIVH7w7EhZmkVSRJkvBgefYbeCPoUHp3t
vywzl1BCAyUaOgRSV/VPW5Eo+p5BMQTUC5wzFPG4uUqyH+nC0HAiow8Ll/rc0JuchvOSDTt38TGP
s5YEikVh2sXbFUex6LpN6EzVu6VOH8Le57Y+3mfSXiPETIV8URdk/INMlcgW2H5HWC1w8GgGv1Z3
YVlkTtYDz/W8LkC+H/7ivBqz65IfKF0fwnbcJEhkr9nQVIWsAJhMHdZR1B0L4yJSBwGsKXAzE9cn
KMDJZmZGDP5xyGgh/gLv6yYinoewNR9Eln7ZG/wW7NeU2+1suLyNHgfN708Bh1wAuy4j3dlc2T7+
TsK+1XBx0YLdOEXfwkobJaP0/sysYwl2ZgDaSh4IPKoSRhHuHX9Hip3J4TODOqVRY9GTkG4Jfn9d
1X+zSDpUyWsS/gcJUVGuH0KFGo6XVKcSNRPf1uOX1G/UTvOvzByqRC/l1mesxkM9GbcBYzLxSMtC
ijvyvh3qVxDuOqy3VHmqRI9IDqcXEgQ643nHU0znDzG3/d6oL4OC4BGW/KynzkpGHJOxY3D/+GPC
u5ixRWbHtbtum1KE800C0SWu+61ucFSgYDEHJwav2AL9PGScySrXQduAeUVa48zrwi2GoBiTu6c5
/kSk+PogQj9Zowa+CCjQPPMH6Mug3Me3tkihm94+nQWoAXB8QxaKFkNHRehp+iX4mjqpTcyVSVgv
iYAfQYTpqn145uvGRi/155fnKRwF0vIjaXNqnFIgsxb6KSZw5Hq+9iWeRTARLVuhIKpdIBgW2hAN
HI1tzWeOJRdWvqhXqNp+UAnJab0R4HlnHM/5MHXOMwQFkJp+oENiC5I67GMDgZukfZs5b5n9uYP5
5VQSkQA4528VS7nsw6ZdHiUTYA52RWdyriaY2+i4xFS97gRo7k+tAZnSyJs12pQ/o7cXk1Mmj8+L
l5/3Et+IPxykIU4gS8BUMvPFYO1sCBcgwX4WtW/8qQjNNf7nOMdzXBtGgcYsL3Iw4+aQNrd8DqoQ
iPK1upAO3FDaYuk41HQToGeGCCH3zlE3Bn6s7CwZv6DjqHdaCE5jivae4gA43cOBE7DdsMR/89NB
lKpkOddx26/zKobnxWbmpBv+R9z0wooNFOEKqxGC8k/6rdc6Jt/fmOyVYruXl8O4Fs8mI1fFtKs6
LTE9ekuH9zC21qQAHGPw1WPPHti1eCTH5/1Mgz1Vhi17Y2yEWhneZE73Uv3+3M7HlpGHKqeyoQX9
Kqt7bGE47g2z5Qw10PI60Jq155wrKr/Fz2oMOqAsG16r60pgH+4Y9+iLcWpHKXdr9u1kgSH3/eGY
CKnC2ENI/CPEFrXc/GcYd+C+qYrlsAM0ViIR7F7GR9VQwy2zzWDc60nTiLS1A4znSPUwcg655Wa/
HMkEL/nQt4d4WqY7EApiF8oG1oEUwxUFvTDKOEw46vNXIUXtSn3GP3DiucLKBiWUgx54nnz4iWUx
ezUL1pM+SkWW5MgI8dJvjw292pAeHfi58f+8q/6eXAizsk8ZOwSdypjEPB5OFCG0J4WY8COOt6s3
UgKTy9DXKDC5wD6z7pFSUI0pIlf+1ZAPB5zpYVnkMP9bnL3RjJkUDE/hj0DvMEtZArqIVndBT4Rb
pnjBVHNaWQio72q0j96lf7/Z722XwaulwUOwiiFIICCt0iVVnGXHPbQkXG39chOuGqbJxLyJ4ek5
nZjCLxPcItUnuz0QsSguIpeBuq0qD0nb45Sb9X9CqW607EQjWBxsSXCkUfHie/WsgvswLLT0kMxW
fnoV6+h8t4wfFsl9yCKJaPJ1ya1wcaNMGHpv12btEdQOWy5OF1vBdJQxDDile3MDjVLaELA0rZpX
Ds+MNU/Af554cqeuT5xuABAiXqsg6vl6dtrJ5fbMtNkaGcT9fi7hGzUkgssDYXdi+iHL1mVx0osR
e4YILYVZWMOQ/O8Tcf0CXOaraWIt6Nd1QMgqanIziWjrqRKYjGlQ6t+9oe2RZmhqudLIOtmjqgHi
HttDaEOVOF9aJfVdTU64JU2zKeL1zStG4lbMS7O/+1211RShJvu3m8kxlYUmMqHKpA+bck7z9hn+
R51Ge9TtZ8jnfdw6P49dLpLUOBjnJXVTy2kYN5AyRXb5cQhxz1DhJ0xcMsv6803LCuHFActkLM06
fU2FrVlQKR4dEU0tEvLieFcIQPCa8KBuBq84jLfqXSaB4kXX8guVMPe4AWqPyKgqa6UdbqmhfKkj
VTlpVEY9quTuvea3jImYyK93hxAL3EmFzz2fjU/PrVM0XPB5fFNlWq8yKI0C8p1E+khYXlQxCQQ8
fhzujnyhcJaAcRuFVaaND3ZvpdY7ilBkcIhIsFmaHXtT2n41tGZnbATfyWj397ubelEBuuOLon1/
bZPbAg0Pb5kzNzAOCRTVN8SV2AqlaDQfbBszgHzLt93K74Kry9ZkxvbKagpmYpVDtk3NCOkbXroV
euJPSY4wQnOL9M8uzEBUjeRQKrVIvyAXxef8CXtXP12+Hj/rF6OBMVAAOH8O6FfRvggxIkSe4UGo
/uUXEFQCpBP2Mp8kzSthhpJOzdvRo4JHHTWdXrvz0YLruyLXAX7qDbpfQuxcam8G3GvSt918DH8U
07G05gAuY2/9BbDahi0nh+SGJV8FDpBhev/fnvfuaoxmCC8atPOC5h7FtEUnaZcYwHXAoSP0FaGi
G++XoyZDFmzAt/qNBgX4hkc8TYLH0HTM4QFPzbFWCzui89Y5fRkasbGNLEM0wm6zPBSsADnFV9L7
gFGFLp7a4Kdd69U9IjSRnlIGcP2XTPhheZcEI7OTmvvqj13UT8CvmXWM5hdJGxIKcx4VjIY8fR+j
YTtnAbZ3tfF5u9fF+6Yi+TtOXqho7VlO/+FUFYZPfqDGSKA/YwijTPHVbMwRQycz43w0QSq6b+Sc
EcEMiR7iRoibt+FUQhI53C+j1IwZKNmfuiwB/OBCUS8n8i5CdGdk3nqCVhp/PHu8aUj9iIZ9c1KB
oc8eN3uj5Qnsf0yQcgtG7rYX9IzadI1cKS0maSOO7ixxgCVVFcMklJ2Zfg/kAUFO6RubguXF879b
TXUTIwgc3Xcs1OAWqY7HW2r77NZd/q+fzK5EatHB488OuuXpQQP/k9lIedoTRHxgIaybmA6ukFyj
wUOImpd+cnvl759Gsh77Vw6F3c5dhS74tUiOybLnQsgrSSGz3pV54rfJqoaXkhcFbMhIW7OvvGqr
6opKzyNVrC5nXCodnIiFEccOd128LfQgsZudtmAi+pcTGNFj8GdT5WjXsJp9Ys/TRFFRlnKf8Gmk
9teWuZv/zPS2waJRPewJOzi/Yzn3gDHvP378y1c7I8tuciqyagOA7XlcAUCger2ex621wIOvKWOE
sB5cKMDg0iYsAcNlmc4ZnQz+4yqOyKnrunWIfxNOggez+90vGhNwrEYAd2ST0tGnIvH3Niw94E3E
UHeO2h/Wzb7FuAwwKfBcCNIzirN6j3vGJtp17QkVqsj0nsSawJxluscK2R5ZAn/guPXO5oO/23e7
oosIXoFNoEGWICrOlsTg9jrXVjqzCZGAPZRGIORVUVnQ3S4FFxV2X+K3P3PID+YPruE5H6HH682i
LALxp72wnY606D+q268mivK8UQTXOiv+TnTvBheeVCnahB69QGRvc62RoWEtOd1HbDOVGHmemeu2
mMYeVmi2zI+ArJBVKHAW1hgjR1c2RzIr+B9uL7KnZ1uktSU7VvexDOW8ONhkvArpHa9wFHx6tinA
vlFcZrIm+poy24CjpzFbvRjpImXQtDsuNL97gWPTyT8Ald1Rmo/1IYSbdB5JFw97rossnPmgc1+F
mg3ojLYv7g/WlAQOKxb3du7XkhXGSKeDeV0QdaApqhdyPyABlDpYa1LsHhUmyd/puieO8H3q7PgB
qnxT7l03pMqPdVR6ILjNSJZCWKvaAr6SIoJEb+XccYLidN6U9sb5pohhN2S2oCoiukPXNrg4vy5t
tpHG86lCSBy82LcCOExTb9kHFvAWTsd8hFxg6IwuvkJ9xoJUsLKZto1zzus3T9t56zPMgGQWJtGc
jsG4ToOm6D6oHXSNTsFSH+ZjKFDwQ2LgVXMLzwmUdLgSvCPJWKFtuxzZctGeulkepQzhFqo/+vE3
adkSxHdDASvNsRFjC/kI8R2rNxRUMe6Ki1GZNWO8V1LPRXV3Z+g/gWSwMCBVxGOdVwmSl5NKThdG
Ri30YDodU7kEXC2Nho8xABsc7tRQ1l7Ze7HwTnwLnq1eRhKxgshn7cfL4C2H/ZNaMJZxlnZ2C2wy
elI4W3LVZ1iXReN4vD2oBAdg0C+TRRo16IiaShqit5+oZDWDnciv7/owNZ0onxHPBYcS68a6ie9V
ZDthq+eWygsTRdu6TOAxxVFZY4EOxulflUMZb8YK9sznYBDmKJvMEmaVwYiqPhVQFSMX8R1J3Yze
ELXwPLq7Zv91gKA1Bj79fLNF8i2w7XdB9QZE9CgbjrZXnTTiar4wfEWlJ1k+iOxNB8FWMc66v11f
y9ypPPvihJ8S92Ue9kMofL1G4MA06j972rAJT30Jx0QALITztMjZDi7PvdI7Q3Ovaq74r6br+DhN
4FLN2saEy8qHw9ggyGuki/B4fja7uH3/MSx8LiwFqP5C+W1Y+QgYS1gKLRkyIREFLO5eivaddppE
qm1AcpgmxGeeHvQ6gBM8zvNSCuIHjS0hM64viGoDLd2VduepkxeqVQNaFN4Riz4aXqAQSWZQhkE+
WmVDkNpswhbsOmGQgL3A1MMaQt2gVjtv9Zoqreav9Spm1mj64WX4cLh+7JL5Su0EWOtFR6KpMyp2
GJVEAFB+CGIYSUnS+ZkIIGKAbaCGMXqFzhudAgKrEp/X7/bQBHwZIh/6yqJjZPYd7UGxDpzgfoNY
RsCjf+5CeblbyBYpRTzt3EUapxU41B4uQ4BhAIzY6sredy10MkEUAs+cv3CUORLhiKErTXTRoXmu
+U7h7fRooEx9iLrUWNUy8wBgrIUHJIMOBcTpxmesqWvjJG5FP1QDOpA9ZVAL2RfWHZa3yB2pV+8R
eSW0ms9yCtiwzSFuEYXGwcctFu2mRsJNZefVQEcb1dBhHojnuoJTrRA8pSpcOCpQDIP2ShnbYW+6
v5gTGkojPM/1y/DM3s2ZP3VvTgKAJEuKYFJJugeBvIE//dfn6Ifu4ndE8QktPeQmWmO+rJiOP9bS
0H9DoctlY+89ZaO7fvzxj+NV9hHJ9lP19fc6RGZuJT1gnUnw7I4nSfZWvAmlifiiVVKn2rduVOv5
LcqMopwSRe9r/58a874uLD18LGP7AkVVwi4BydeXTPg91kaGCcYXo8sudUW3o2eW2FkPdGVHZeBE
k6HhFxssyhUdABXjuzrGCPsRnqUKzm++RgyidnlkvkgA2MXa8akHqaJxQtBSVatbUdBuuFvjEbwo
nrapjwOB894Q6Qw7fikTA1MCwm9QkXKztFkZoxnpXb8cz96/iTn1vKico/RNEtXQ2/Xzq3NfuW/P
Fre+wR1fRotCBmwWs1klX7AgupSHSeYcO4pLF+C/HXk03MQBTsL4imhU28v6f/+zCkqeOnRz8vqu
+qucXDn8IFLtkQ1hgc2t3sXgDAQCgIm7Y+FktUiDPgRyIM8bPEUfSTeh3jprbCoeBrDJNdtmILmb
SgaANmKlEIpeB8wJqohD+JuutKzXS/IjybS0zvs5fpQq+weipJ+0DshnLOrl+9olqLKOkkgEnRgp
osdZeDoKpOylqMM2PoxDkJLWFGa7esXj0XW+tId9li3QtSp0FCV8Qltw/+dyZagRFN7UYVFWJpF7
LHEI3tkcKgyT9G5e0hr37WI9vUCFLGryIkuiilIFsgATk3SPomQp/OypoTfBAviJPtNwsRtHYNWD
8dwBq7RV6/nQdyRTk4EJxoTvPTpHpf9l0vjM3ZUjjCifOKTDU7zLFR5+BhoeoUbKLAm8540QSxI6
f/eiFXdK1/e5mZaETWhseka0zM9rPUGVBgaKxDYz/t6xeuPVTEr30jp0G+dQY3qZrLDaPUTNtuMb
Ofm3s6a4ADH9EMr2ixBT1QHmGxUnmIc3d8h74x6w2w/3D9z4fc88fBHXnfIccDstMlucHmDNZXtB
tGvGhwLjZIttyukZmnDetIU9EeYT78swydLyTqgCGVC2gQyTNqWmAx+3t+AvPVuB0X+q3aEoeDt9
HwaT1/pqYLVE+Cphi1di3v7dHrQmlZ5qSuK0pWzVrZKm4PEUYyOJJIexKnacGTsWWS1kXvcss03i
BI+C/EsLa3YrIJ1Td0g+5l/1GYFCJJTZYGTxQRL2rOpcstTRRY+q98F+IKt1QiBwhYiLyEEf2t6D
cCQkfKjAXx+EydK/KQUyhenJ//IZxvOkCogSteXs7Q2Tnzcjuw22MPq6bevn6kUH7HyWXYY2WbZ3
PtJKcf0zinZ1LiPGsOiI0rp6vq1FaVIHU5jl/eBpdvN9IyXLAHz500iZCTlULYCVVB3wial6/lCh
0M9seqgHk9e38ycBgZ1nb090rvdW/n+3ksxFN2E3Fg0eibPL5nkwiu8fP49q3VjpQ8j2IKhrJSdC
X5q4lin9pwVcOdDs655bXpSCgk4MHKwaHJ83GT10HqFsyJlHYfyOpavMsPcuQBPjkM3+aO5RVozK
mKcNbdWao7RTkBHq6eJXb8A7N6JWVaf4jxU2afyomRtZ4JNxr5UBntiPjyBM7coYiwuVnEzDO2mR
ISibl9h+1UrmHMRC1N1N8tJSUQh227jbdGc922kcvFG0fEev9LfadCJdwwi4PrGd/pXlWhxdIQ4R
UeKoklqu+eXOCsJ6UWi3a1G6ShDdPBFqHZC0NbVp5u/KYgWi/Iafq00QXybp7/+7U4fH18/Vzd+L
PYX50JVwTdVBmSngKJnkVtjVVFsnG+T9+vDKWkreqhGH4DP4wrqCEjKCsgHm/5VUryr9Yt4IML46
3Hspl5z2rhnogVtzLKvPArsUxCqk9fFloUKMzBQcem+XIQ+H3LXDrcHXWYa8pt5OWANm6Tyiq3zK
dKi9MKkp+ckHRURMWr0POqwAzEnhKB94pZ/XgxPGD3wGm42yagerhvztheuDYoFv94Qn2Yso9qhE
Lx3s3HQgqWrDq9DSL5Iafpc3RuI7I2bX40+p5X+d/AbbJMzLu2hoOgLw7Yy8eSdFOxzjMLM2Vop5
YEHnhRKLKOcQcD5tI2wpjK/DofnnFurxWhaDCFLyMAVARMWoYXrvbxiyd0yvXrQjKRw9c2uQyTRM
p+BxYuM1egc3FbBSto6vCPhr4E2DzOrfmWYAlO4R9jOVN1n4irleR/X4SdEewMiIvaQuuKes8GlS
7idP3kFggE6QcBjxgyTfFXB7G3iXWV+3JqC9MJY7VqD9bWfDHc8Z+Tk9I7+SQe8Jxsyt8Nt9cQUV
AYH2sTvQSZHajucWiCGtqlZIXafYXzDxFYHQ/Z4exjXSAVhnIxElRdvz/AVqrCkRmfdS3kJ4zWwr
fOtsgiD61YnwVV3HNF8Qt+3EoPcnMo1HHdQOateCGW7P2OhVbcWHFX2qjMXshukbWgem+P/yWoxc
eMnP9TGwq0wbOVTmnxOMbUZZYYQdPijmysDh5KZoRSY+LTdng3G7VLHR3MK6DfvqShsSvWZzlGB+
G+zWK/I/VodHrktQuE4Bw6u7/wjC4AN4SNZyuzApnzIjvEF/smjJGT8rx0G7lmPxlScsdFwvfL7j
gGOQnO1VdMPR2heGfieokAnNLLatalbYJA7YYC0+oZsX3UKADXLRoX2IhQ6X9WoyKEew3kA9F9Jo
7iNds+mHyPZQai902QdZQXj57qDmuEhNH4D9FHXLKtylwBeKh0xJfNupNwMvqQytUcpUoPZnCPCt
PyJTWnHs98JqKonbcjhrN1cZtY9iSkf0TW/fVTJDaQKHOgyajFiYBYd4AL284O5jtaIsYQldbZQP
2QYMObEXZ5NvtA2fqRzT2IqPekB+eswZzGUIpYrZz986giR7jlD9cLE8aSXGaCnJf0vAPEIKdAI/
Tfb1svNEKMvZliO6+B+rEUj2ESXb8kuf7hqhyO8OdoZyH/HjVO1njwBQE8pavkm+CTVeZVj3FjhI
VGNRlcw4p5N4EuftOi+fQI/PsAL/9jv/vQOVIA8kDIViz0LjccQOnkE388P387d8CDCwGXc8i9sK
BuGlWnBx/lhqluDwIxSt2jU7RcCSxV2BcGB2GwrmaltMl6Q5N/aFA6PXx4fVojTx89Xw0Q9oVPAw
Ji9746IshTAUpiUHRMYCYq+9YFxj38LCiia6eZzrPjk3OtuUR/gXwk9+CLzc2q2zmiqEffhDAaCa
BJsJIbjMnXl0nBHHJYBUr4j5D77A+2IE0iFtSnm5/6Hq93sk9vftwyw1RxVLus5cDLWn33uGZMWO
YgHptIi9bIuqYkEN9Pw4ae6xjeZbahBpCm2MNvyrZihBRx71dTRQstuzC79iReUkADQWuCZfwG5K
8myOzYU60mJjWGfDUXkkGMLBXkFfGqnGVguuuCIEvzScMV6ypxkhq5+l1U3SB4Bo1QAzAmaPMkrm
fTiU7Fq6Gh7mqIXWgkj9h8dL6s3s1ewsjyr54PDufx4/dzZKgdKMyqFG9JiXDRIl7mPmSqDMiBmC
M6y8KtgtMVtfu7crmyfHXEIM1kCtQFMlgCJ5i9LHbuF1uxVTvYi6DM1BoNM3D72XjpD3GCPAGUof
PhbCZHCV2N+eFRG10TQhYw0SIX0B+UQjKBhVaLLRVPS4VTkHjM8TJuGQpI7mIICew1nLBiQTCISW
vRWlT8Q3As/Da2FZSq9fLI5Rlao2exw7QP7i5vaFyhKVFr3wchgjElmhZJQiCwFbTdrP3E+FNtvb
3AiJuuth6WxlFINzY/gNnuZ7P42qGgpIGDbRCjpaqXshq7KX+zbl8s8+FNxt543zbPaqM6BGvIEC
ohhymCju8xsBu0kf7AcvauinsrcI+VkGAHrj7iD9DnUCjB3NtW32/RPsCRrRbTrWEOg4yLA5qM/V
ayZsKrTdLQMptRtQCLyEeuXfx0c26GLoHW0UsdiFqO3+jVOGuoFZadVdNcCncJaSIDXHfgjMO30N
98ijeZ2Pd7CkU1DUAbjPPPFEx7awDF2qck0+n4UyhPx5slj6F7YkmelSXfq5eoVwXbkWYGNfXB7G
IAjEd1UoMnKWYHbntikxPYJNiLrM7+7aisYXL2ALr07julea2jbmEsQYsBXCVZh7EUj0w4SjYCPK
XRolrO/y7YHh8gi3Lz55Fnhs/lsuIM7yJcsRSIvwPv1UYDYVsAZFMG3DY88rcojNPGcU3lIHQsgY
1N417ZeEL5bzmoiWwxpY/CSOL9PfmKYolB8Xdj46Nnm6CWYu07bf3Z4jpgMzdpyKfigpqP9h65GF
kZQ4iDl1GvYCZoj/5lhodMz/JMwotApJ7act1qcZsd5iXFDS6mv3BhgtX1HTZiMwROmm+mB4C0nc
BSfH3rtBrzyrbRrGcXe7EMXFVxR3EluF2Ou9lf74kNajosJHg48xvU1C9JvTXg9Gy1z1nbAwchTE
tuZOcxyr4BuuFIhc7mw2nzG39a02+Da568nv5DdFoh9DdxWbSWKNYP6NJZ3NdQSj8t687u23lwhv
6+DsZM5+aXmXoUDuB6FKj76vCTqFuaAVi7rDJMNALE9zcgn2h8yGZu8NneI1DA1fYWeNIY0QRkVi
cP4wPoHR69eAH+zX81FD47RXh3PKZJ1SDgvIVu8IkeQK3q1C2ECIN72yyi4aV/zEsYuAvQRlI9uC
WbCGqe1llHNThEOZNyTTF3QW6PXInGVg1rW11xZaJsCobs6X6874jDC+ti1en4USt5tMpfw4coHG
fZnctwhTsbOda6R5SKrF9tvsHM3GLadtrsiNkNoasVGY69V0B1BuajpjdbB/fUKumc33ycURaH8u
zZTS0HHbW1dzR/NuRMmsFqb7RKWLN7g6IHDwLW6sNTdMRlEiCA8wIvPQR2jTTlWP3FJGThTbQxvF
bowR9Z6MUY7f7+/CBkLYTudb9AFJJSZaRf41xkohDn3MoNTE3njOQNDfrJNWGpYzrabPQmztuAK5
9ICowIyhjA/ss/hk04pPXS9zsnr3Fxeal/oUblET+TYwWQ0BM2mb6s7OeV1ktDsDeNnBO/QkAYtQ
Gp8rCywTHTaOXsnOPuqD5Z2qvwGY1WZSNdHwSzgBX8GO9jBYIfkLo/m+q9laN4qGXRM93T/A5tyz
KtLFwvRLdYoV14zqWFLP7PpZtH9xDs1Qi5GkgngKpffM6OVZ0AHDWLj2Gh88xSZYP5GgsYHOXOki
FvIG+vOU8/6dCCsf8ZxC+BQDq51D0DVznpLih8bQI6j4tn2+9SRvILUtS0VUeHIXdFUPG2AywE2x
iq9OEp5m89ySVqlZlzCBCZCqKK4u+9w6YP667ftyAKbZHr1KGf+O+p/ne8z21NUlbFQjRtYt9fnx
wLOqOqQIJItlBycnzbX+MvUNp1wRhDKpqYTd9kJqAm6dWO+NqeptQQHqO+hEoSkkye6FAkqHbizV
9ynHR1mlXIh/JbDznCZM2YkKps9VtLYwo1KBUEbBNeXTd36BzjuIVpxKk+MGf/Uqp6PD/wugqst3
9YazowBgrTvB4ZdHmPM0GG2XBWCBXtnzvSzuKjDtke1WFKua3CgVIVt0PSG/9necVy8gRSaA80eL
uHD7ZE/f4sV4rg4/ZGYSPuQYXmMJYf1fGuFfLp+cofMowPZ8U1ALz7nN2gvo8Hj/BsC8PMiBQt1S
hLqmab+NXqjDgAPND1N7bqtpFgBWoXAyjYEjJcBUkfMrCxb5JkAqhjGMxDDAIVLLLjGljWPvT3Fl
VB2WjpcXke30hPKVRqvMKikRpWJiauaJMf0IwGlmJsOYapTbk8oqvDRo4zBBSTaahJ7uOHeOnqW5
8K/OZwCb1MIN5GiDbURcgG8XJunJp6rA0DR0OserejEKS5E9qckYc7Ru+/rxTF27bw+JEqa2aCnK
tmIDSJzkV3Pba8xX91hDzD+XWT7Rg2PAWUsjS2Wa9omk3hy3uX+VZB8J1xp2wKi/YsHGJB4u7gdw
YgNeolgsDjyqC4cYDRQRqJX5qn8koqTk/Gi5OImbjOnNPwHqd8pw8x983fP4ufhEX74OhuflQe/o
BtsBEoVo0+Y+x+8lLyE1V4tQzQAJyRc0ed/VF0ChKJrurao+Sr+KYZttqC9c59y74J0NDvx8Yu01
ghDbVQUlZY8j1kMndjigVrfikHj0oUziKIURCE/hw/9uGFqHdyLB0vtR2HvL/CrDOQiwrsxdcRfI
i2AIKRGCbFrdtxiHxIX72oiu9tjMyG6mtaI+lR+d1Rv1THsutDVMjruSopSktR51z7hU0CzHatiY
2JsUfpmI7d/k4RWS/fyP63hg7YmkXUS2RRqOIUERDJm5hkagR+UI4iL5aui6d4IkXsatbELV0xQY
wI+JQvodU5Vm85fVO9da4VEeGlShaSRKsy2Mqugw1dybPCRNyQnVM1QuhgnEI6qbqbeKrEhxAFOR
BR9oj2XVME0QRWIAqscc6Q1npHiN40WDCEOqNopU3hSK9anjUhVzFRX970WIv+GrtsM+PLV2b6yH
7R5HyAmfq8FUVaynKuwb4P/kKE1kB7MjwZETyKqLJyRG2fZYEgauwiXGcXxfXnI+SViJ8h72j9DB
U2C5zIXmryLqeMcAyEpmb155T5+u8RdFLlY994H28yv4CuXdTq52XghnXnvn9x0co1kMiX3u/e3N
pPIVjbtKYUkXRWIWszbmeXYPQZZTseczpy2CzQY8F6OV7gHoOL+pLkye88VW5bb1G1iKkfpb+yu9
XZ+PTFMgGleBtNrzpZXJ85X19koG130Qjs6VneQ5sKaI2OkcUJsEn/is7Jmwb2qOIMgSujEZbpEq
AG2+ddqxXDdQZnoiQ4Q9s5fnwsovUvqdONyyqXvUwmMoMMVnkZ6FGJEScyZp8Ycht7M7MYjsTz/6
WHFX8vKe0MIR1FxbSqX38HfjdKZyip6FsEvgOsJPz0bKmTyGqOI8RY3Ea54wQkOl1ktRMbdGU+rQ
j+7WFlhbO1Ng+2749x7lthuK8aF1L2TYjEZ8pTgMUc1m11zOj4i3kLNknn6b4a/8NtD6UFB5UTD8
eqf179Y9YlnxfasQPMRlJPF6lHjMXokM5jXHhDDh7F37kAr8ec3b88PwE+5sE6XoUuaWBcFAYEYd
GEJvB8yYUb1QYjyOapKt/VEEq6/PqeZT6HS42Y2JrwSAMHlQo8MiB4o4CMxN57MXtfP6kI7p842s
ZgbW9r8FKshc6PTjcEzmqHaaFMGDq8IVyHeDlDf0vaCFLm7RE2ojL4K41Z41FzQJYZXFHjialciN
5wfgotoRgwYHX9sjpOQlbA3J/cMuY8Krz5C74J9bqQX8/zXSWFUBpHJfeXegIwmJw8q8uJx31Wpr
Jp78IPKgvb4UDWa2begVwGRXG9R+dMiQQj9sxRN49M44STp9Hi12ohIG2Df5b+ZbMQQoJP1W0Tnp
dJ/YI+kXlEVuoIqDIO2NN/Ve2KE8f2w7/ZI6eGNRjyvxKJsyrL0Un6XgRVPzsXZZ154/FKhQH4T+
rpRp4puj82UusaPd8+bbL+Od0r2fclwQ71GXBM9E7KM/+QJLSzl41ySvNB73DeCSVGvwuTRxrcW6
9Fp8LkoFE8T3VMDB7RM8WS2K0ufW7lHxQzItFzVTCTllr+n5ZyCi5C5IWmdyhiXIX+QDVpzVod+b
W0rCRIraiNYxvmE56ENAzCIb9vOALrJtC/R+SH3nH5QfsYjL3g/bIG70CHRdER/rEmTJAPQtGkXF
hHxmmMvtCRt8cZFrUoWIDf7BMDDxfnCy0m05MS+OsuwzzresapdX4RbfXzuYtDtMrIgK86D4aP+A
vQLTuSqQywkwQzh2PQtMVoU5xkmeg8mWHzoY5440p1PirMu+Q7yMDkYcNpeudornp5TmiaBAXAa5
TmM99g29l8hvvLGOIrByL+G0od8rQzKkPsG2KCg04AOeb6p7urA980m8Y3lCXiZ1P5ODN8x2FIWA
hWdm8uwyvmasLgiyThw3D9Fa7bxkUZqfjFIWmEdyEGKOb0hrxNVp7ESZtSASEnFignCjsSGu5SsH
ij6wY3Uiu2/qw2PQaeSWJWmX0M50sNYBFWdhYjJHXw42x3/CDWlk4/7PJblfOw2IErEGLx+Ga+b9
G0WgQK0njppHPAmWNQGiSu/6NsKFuLnEqtjp+SvSdQQHkw64K9V7KtcTcDN2t+xiz0fumiuoUbvO
PKTR3aCSy5MR1ofbRrQ+1hEp+3bifw5crPuZm5LPeZC/Z+5EJyoIOspbLocY2byjo0/HYTOM3S2D
ucWgmG564nAKGPE38LXvUUYE1AqHXofR1LGyp4xcQzJJfnAc0aJsiG3fQ3e1pRiq2Z5ImM8xyq3q
MPqKbin3VyMCIbqEkkN+BbzU9TSMkD+O1Mnte8CkSatBQRQEQ4/NEz60BXszIm3cnmLJnnVVaVf3
VLbQRXH3nC9g1ZcNZ+XEgSeXHjUI3Z6+UFanBAt9q/BbOKzkxzZQO0Jih3kuOjyO67MdHS4+aVAY
6jqJLHWZz6TbJZ1k0Dx/2k9qmGBDnHJGeZo6l3gzvI7ibXNkm2Gi7rCt7GuCjaWmtCe9Syzf3Bhm
VUP6gGCVCYCuqd7iCXvL0DqTRe3G/mjEqTVIjcHUXilalZ3M+MO40unMfabHhv9jhTE3f3oiGJ9r
4400yAPrmwg1xHwVFGSASJZVVv/B2JCpVWbjcb1618FhlgQjlK5NQ9j9m5Yzrl5v38dxEqBsNSUp
Yg2owt3jv2Sv40a0kGgc6+Nyzc+n4FUruCtEVNGrQmVNqzuQGw1hlWIrvpK79ZlvdwSxqzPiBCGI
JU/RxkrD5iXrkb8BSGs60OhHIePkx0OrcZPqH7KoVhovVBtW7YsA5CyypUitY9m7k3MhPQ1MFujW
yRGaKS1WVPjUoscZm7Sw2ER7cm0ru10Ldd5bgoUKvLE/08rFrk+ilo/ipWW8xzP6/SFgxUXmbVCU
874D+BSsGlD/2o9nzPwwX8pLw7Tlv0NP+RuMmdB32gWnfTkiRriiBlK1ZAPkxggjx3fomcp+CSIa
MnV0CmHJcnyHahJvA+leKWqWibmstukYp9m1M4UMC0NpALvSlT7tAgHxVlvL5AS1UJa3yqe8YIAK
D+9BxFAGnQKCIsvpvC728KUbcQq1ovpxqw0YILuzRLRrmpMS78oVOT9Nruu6E8svEgP4hadp1/Y+
w5IxadxfXVACxyK2WQDCPBH1SYC6+jGfdXX6GoicDOYfHEaJC3wefWO8XkWjFtey6mW4Ql3tqAOm
nz7J7ZdW9ez2xM2/D9TkB4zah3x6Ul7uFwSQKFdMsmQjFF9nHYqcAgUaJux77O/8a8Yf9GOVymXD
cmgMfOUrjyVtzEeKUAgf5Lc8/J0bceNtbVlpHiNx6PBDESmJGfgT2kPvsTaf1zF9uaOkTw2Kjmv2
0GXLssCTi5ZzdwO4GaRzoJmdKOdaDFML3IyQaBMusyRcQlXSFKsHusZyLiAEw5DmQggY0W2sZk5f
ZjQ1lCI3Y5C+6iHdDiNtkiYsxlQZ1rlaNsXSd6O0FZuw7jBDVxxTu04cUu7h1TD1+wAeRVVuEw8s
/0/7B5rvYnvqq3npXOn8lIeI3JhqX/rJ542tlXiPPTFadMEK35DTBNRE3jC5WANNAFWOSu8PWQAD
cZAsv9WqCiGJctup8BGXq3g+g2nq/+WQvRzWOj0hrn/a0DXu5ZN1l2gyiktTQXaL5oGF2+Ymx/92
Ti4K2BpM0sL1YkCRoCxRFYSeqUeXoF1T44SKX12txCtY4rzK4VUn7p1f+dZEJVFZWLQ2XmCbEtL+
VA0hFrLO8Qaw/CUOha90k5nRRtRgntttcgZUrU/TqTwiZpIzISVIsUD+74pIgCtBayp/sye3e0j5
Qjpdm/dU5rXnYI20n1G/pwCUDj1+kBiK3jI97GH9HyHqjt5yfRG5mniG1kp2iboLEiTfbCu2w6zV
03KhWDKt756H5p2VeJhJk/F4bj0eQZz24eCeJh6C3H6SWCmx0L0JTCalMR1KZVCFoQgIo2C9tMc3
PKQumVYgL58zDm3IfIuwgQYVWNAa5Dzvbs0PIJxQa+H9/+pwfv3y6RzSuUdUSl/cP5jvRf4BcK4d
ssvadvusY2hx9yua2FKh4De7GvH7sYkGfOk8YECe4FUiyfdp0lHvB2+P+QLHk2PetQhU2l6kFECO
xzdcsJ72lI+uEOtIT3dUcrtFjEYefP/INjIYqBp3U7VU3YTGyOz7aNZmGdDVehGY1dOnEn3fAVlp
BH8X6SoCKGaQL5LVAXOHHWrFQPZZhYr+457XV/7tWk5wa1HxFL0AKKDxchZgp01Mxtfp1bAmnduC
NCQXo83pZT/0d07kMQ4gqPlK9Z2bWHLOva+ZIL62+V2KH7vSTXG66rjOOLDhFwQ6Gq9RO1J7Tmwr
BK+NJQ7gHRmpqwm0YqIcacusDVyMgSvXHgeOfjwprxiqajgFw0BNYbNeywIcJatn4c68inWDHaHF
NpwhmyCHPEJIU9+ZmB8nwuBxVdNkP+XT6Ul5c7sKCDeF5rpip2iBKVzIGey+lUKuyI9jRGjUIYkj
FqYpa24fLU1tgXIBNxEUbkH11TZWvPltgnhIMql8mBnckYjazhxI8fhwZ7k+0YVxshTatxU6ZAHk
Q8oI7pUz7zPmYIBNtP/mZbZm0Y3fqZdbOv5L269Chq/fYGNa/SR/Hw3kCP69q8aNJZdNOh4U7as9
iwK4/ljDyaEvnjPwdaRdO31AkVh2q87GSVfZH8q6sW4T4dFaHtXnD8KtATRVPh6k1NlNeFSo/hsb
X4Nh1/lF5J4lQsXPsUi4wJ8TpTfTui0bmSR6XSiNjYV7I9VXTF56rmJ5L7Ms2Kl2CIfQYFhECNf4
9jszeDNv4AhHiXz32Jc7FlM3FXP1A3aMX8UaFhUUL/vEPwm9JuPbx6zb6JXu1Ya1FusWyamrnQT7
AeWRRORdOPEiohvHW+956clI6sFGeelR4KJQ5/ha0GgJCPDLDZF4gJbbpFYGZrQS3dSzcvucIkYo
LlC5KJ39EsNmm6xuGxnFhpfMe1AcSH1T8/DElQb0KGuzja4rcBkQN7lA4MAGZczVXtcskvuHG++p
wMI3vZm45yvCSiBLZY7WDFbp5Gs+aJ9uMvyCtpS1AhapmKT4yPv+koOuP2pDkKE8bMsrmrd745cA
gsgMu87VKfvysZvMRTmnINg2ovXeNOxMI/v+NAjHDYjpDjHH3pBimUCw9MSAl6bUSGMyUTVyYR5R
4ot+X6PPT52qD4oAJ+MEljYFN5pVhRFVqIfPnO18KrDcnTgIN/OF4owLG7bRjKqwDBwz92YoiGzj
zbLZBPXKkNyqebG2kvZR2hZwWgyL8zL45EHk0xvjirCweTxodEN+UMnBbNw5x71pi7wgy1UxZOI5
a3VOEfZ6BfPeb6cuY8ari5w5QoF1Xs7k2PC6F7ilwZ8gIlUp1FR1X9Xc7jbkyiypXL0gfpmZppx7
3oiMZtPzHOwJXrCrTsVxeDaAGMNfVe1W1UIYwCr1/KplGzi763CrCTQIChM3gymSBCykUQmiY19u
tfRy15muaw5vzEUS2O1KdUo/DURr9B+KCnqzb5TdfguMqUaN4higB+59E28xoFmhTaa63FKbBim4
swNc/vNsmvXzhXkOzg5+HeFddaZk64bVLi8zFcES3x/Sh2sPeZdNc4zEVZbot6Y0kjWBWjuhk+6M
AcJWt02Sc8bmEJE45YJ9un+Pp8TWxm1CHo9zbFlEO3ZawEbZzkU5NMLU12PFhPonVOQu1ALMK6N+
L4IU7RB0AWIkXJemgiFtBIb9y0FSp3IYnPssENDe6GhNadROViQ4CFlcGlgFgDxbkTtF7UUsBq7f
xrvezg7mQIIQqCkYEg+dDhXkGJqGihBFxvnmTWgo71vB4Uka7GQyKIo+7T6EEgVJosQ5qhioB2RZ
ih0Lv9y4qfgwk31v3QjdvjyV6s3w2zCFRWOrpcgtcezUj+Ym+VuDxxEji4RjPEqu85QyVxuyD46c
wVer3WSD+1/vg4dCQl2riaIklQyLhu2gf/jED3C+0XsjCkpX/99Ey2Sby/5bWw0ckwdvqqpojxFA
7pyMiDS+nFIsPaZ2AjpSVPyIrWdg8jEcsLa1psdxEW8wmzbEyx/H97ilOFiuM0GZ4AE52NScg7N9
U2+7GVAx+cmy8kyJXou5oibGWwPgA88tyX7GmIt00zTycglT8f1qyciQH4yTY+rM52ydhN1FShXd
/mRSfwZy0vcMyQBUMktFtn926xElAMIZ9kFbcUaLamq8/KB6kVpo7YMxHpX/syRj0YgKHD8ArngO
t8sSGz1qHTEGK0N81rYpdzi58JLs2a6aD5JwHkDdnlibh7xEIJ4VKVIVqpxCi4edTV6JaCV7xvMS
9Yaowh8rUZkoy6z+wIoTaL+FN6jMmQfbMctNUWgKrdb114ct8oGkMNi5dYcD/xeWVmMEMmTbZM2Y
AWByXJPMyQrS+qHGIextIhFZjFRzbVKdczrYfYmZ9KTkgUjMcK4h3L+UtwvrJEi87IKNMKWPdRol
Mbesr4PM8P8JMLxEzi9UAqYIHaDif4Mis54eiIGBbPPzbphI2MuiuQW70mpmZ1KHqczRWWJYhd1Z
froDWXI4qNJpbbIGHmlJpB/AtRDcSXYfP1b1n6QSboTMgrB1hK2y6vJ/CNt8jZUaaKkmLMC4nyxx
usxWK5BH9YXcDxTVDBNzlcP1QUvZYgleqKkri/kzt8GIFcXMBmnQvEZu9Ir/MdrRmR8i00HEyEE5
Z4ot1gVuYXioT6D9Sx3dL8o1y9OM8xFgdoCAsGVyrZaf3QOClM/e5pn3y/u7UPsAP6u0NPI//AZD
Y1xNeJDjjCAEs8ygF/PWTp6Z9VIA/g36qw7zDyd2LxseCqoclq5nF0InhPTuMvZ3L5zhCQQkgdso
Td9ygAxaMK8Eg+z3aparqQ8ra/JNxSwHkdEbMpYn+2z7Ca8t5MYkDgdd/DIKgbfKBgSsjUuXG9QI
5P7gB64a5DCB9Ovj1BY7gKE0kxriBfr8wigl72J3gh2H+jMvE1X/OC3+tcsDaF399Z54mkjYNFqe
sHtsWENxc6xVXLf6tUK5Dv6DCYcZolEHzZ4CIShMwcHdnC8q2D33H3CyB8IMFtK25mMRchQIXeXD
oYHMlhIYIe1vN8bDGUZPxdKT1vAW19yNEZMkXA6ys6lcfVROWSRXvhxDH4bWwkqw5ySbTvXN3TM0
/rMRoqx/h6GzJU/TuS4N/yEM/eRuZDp3prn8ZuZ6EANTbYX9tjz7BPsDm5578tcrg7aYH0ROb4eu
zQ+ObQt8k5/Rz1rdRdu3XK/p1OplpzMp7cp7mouaiWumvndywv01Cld1+nRBpImqvNf5npMc+ar6
NYFAz3jgatc64a02OOrldohnCPaIDrBruIoXz2krL8LsZZ5pgz5jYhqx5bIGiTjs0CjdkbL3/y0f
2i+PaxTRixp9jV2UpJsDUuLx6BDGP1gbGyjz2/+3ofPeYrioTQ+ll5HQFWoHE5G/rdw7Rlu/Irzh
4ug3NRS4Ci28hrWMuKzcMS2f6pZ0BydZwN/VmLkvchZaft9PDSZpLdPZBVHd6UyvLljtAzmjkl4F
EufF0fWTT/0hsiotL2KnVsx14DxNXbBXrW6LOXvHuUnvQpr7D0j0CnSEbQiyfQFpbq+aWuUsZnyz
zudU23iUMkdAmuxM7w2mWQ5cMY77Tqs6Nop1fdOOQZX5IQ05GdKaKJaTnEqQUR+Oa+fwfUaPK1JA
PtXtlEYONeunEd+WGVYm57mmdhAO2y/aIDWpsZb+4SqjelX1+m1qpLwTGIdsVI1zZ697vDp+QCMi
olUow8dybwomf9JcN6u7DDXkqlQhWsivjo+rXVoK4EJxyueACjsCPcf0oarOKH2CLV+YNdhbGofW
C8fsel3HRCzQsUZqGn6EarBBCoLXjislzkiz9eaa79Qd4w0oIHKK20j7MI1JhJljqfz8ZbB2uN8E
+TAxhuxt1YEk4jeODWHE471spu8pb9v91lHnb/vhjWomAYvXXC2vGXxOiPLZj9GFQyp9VN8tc7sR
zhtGKi1fZw5luti1NHsmsRTVKGOJUtRBYCvF76U4dwKrB+6N0i7Dd18LwL+W2s/LC+1NbqAQgkL8
+UiDjjpp7psceee+C2acjl/yHtu3A/MNV9gKO8X9U4unBg9dSXPE21MYJAtgO/utEFDoN80FHZec
ViSNotGQpbq63eHuiaYfty0rU90GIjPyciMbTATUz8UInamGYA2mYmIKgHRfhjI4Oe37zHXzWDBZ
/hBRrTm4vfmqnY+WEleqvhfLUoICGKPoU7VyWpQqVN8HiI5Ikn43Ydmm2/E8CnyVYa8tqCn+404a
i8bNzDbbzhdbtZsIVwxDpPHe2B0rH8rn8V/3UY2UzZrdW/vc/oJFxcEUA0b+D/TL/bMK+xhQju9z
ldCtJD3xKEEydjhtVArcWuDeb+G94cRgdDRPOae/qx5IwSG/h7FPW1rSOgV/+KJ5ve16kN4pb9OI
cgL7y9a8WxBZyTZIm8vaoSYUIx7vowsV7svcRujQoPqRnvwZm2psZB9/gIyIi+Lr5RwKL6c5LTx+
Toh6rzQgu2ryFPunw77Qo0yflEhM5drWfv7Cd9fAIG/rVX/mRjLkSOrS1aodiD8gqTi0DQ3LzVsa
ajoyLic40vd43QFPkxxNibzsjYX4gsg4JIMM2GVbVbEAssILKwVX3Gwukbe8OagokaZG78NH43nL
NbTlGSUSNdsEAG4HcYwW82OQmcN96j/9DPQvQU7DggnYz7vzcqnru2LSlpWrj8vOaJSBrDtx4niI
XV4glnNU5EnNkXhufSdRFrHqbep16awgqXB0pyYieeOnSOMvZyFPWFwhIQSWOljIl1Qgp/6VJdtB
f0taSb6YNSxkbHu/uwjDo7Tzv9jO8ys30Tsv96j6u2C5fAccPKFYzWXQo1Mwx1YRvMGKn4Iwsk1/
CaJ2U637/675VDviELqnu+ZQriGQEx9QG23Wo+wrYRkj0WOVXLMW03kr+rwmfQWO7qOxaSf7Jo5L
5Zi9F+EEJByvl9FWWVMi4pyh9V3X+CeXhNo8ZD9Fb4lGUwbg7OCMW88BETkms6yY+urC2qLfaZPr
PVhPiHiL5ZlOlDvlgHFTShbY4Icq9tz0RZQuj3Gn0IritSui6jDPTXk5QOFpA2ZHUvRIrzaZQFxG
Xq8pvZylNeQ6F9D1DqkmgOuRkgE9HO7OnA+gHczTlCWfO7oqBfPLEAjllymTSQ2lntWv8LRj5nP1
K1zvla6VnfaApYZclIrbes9NeZfmdX9uwHp1oXtofA0f8KMqT1Hhp8wxp2/NW+yFRchsrUofnXGN
bCxRpD+HJi8RqtStcmk5AvGHvD7NYnaz+UdqjIc8S24DfjeAFtD6FaQC7Pza/Qp/Ksj3A+IqnB7C
IAt3tXaUth1KMpgCOu/RogxCjMO2EPTDdg6k8+ehve0BZL1yNNW1f2kNYqJEIPN3afPHqcJprVbr
ouawcuD47kvd3mPlSVPzr2ZRQiJBknQE7t4fALE425Ky4N+jpdSCV95iYdYgCFPQxWIXHE9hoxUI
gMN06JOFIrLlzCuKV7BMRZVl5qFZAIHvvXlMLMVE8pGZ+o7bedSy4tegEdrOBfyWoCgFkHB4V0Fz
7L+koHtQ1eb5cycvV6MVkGhva6P3l9lk5VNbbpHXf8Nk5HLkCkKNXvWYrFIpH+fduoHz1dQpjeUg
doNUHSlTZxYRPiCYR2JloGeyQrS/FAuTsfQRyXwwVS6Hp7en7fP8DpIIjVXF0BM3RdFAdfaoNcJX
OC5UL8gk8aqGbtHAyEeN4xAqKMvzIHzLB2iu0JkVrECq2XGbytxgjajuQg3YTV1YchXFtkKMaEV/
PwUzVOqEZ9XI59MC2tC0C4XZRlw0WIX2Ng7pbSjJ6t++YyokRh6Uad8ZCzp9i9ePT4HicfK2d5E9
ZsGOGmSQvvvakcCNxSrrxAUMeFG2AYPlpCe9x8/nMWgJxKQloOxX+Pv9bL7BRC9nJ+80Aslx5ISG
WAjgWJYW0XJXEg4KDSQwrh2k2ifiZa/XsLJvVixZ6EbQRIwXWhkhP3cTnE7dFRpOoToeSaMi9wji
OcBSm3ozJuE2TjTDgrddTKISsoYLDQETgdpSwj87LPeD2OnfhQHNKSunX4DBxKG+j2bcfsn/7M5f
KjEnQd8nnwFHUhZH0e1644x/NZObiQHo5GgWnXp5b+E3e9nGq1pjhw7l8qptoI+kX+Ui+rQE7ien
XeaQqxh29acm2djBntU6XjlYBovL9lE+5uVPeocI2LS/kMD/3qaa7qdHQah+eEuXc0TxHOXom6Xv
8vWcgW6V5XiLszqg/tKtftt+bRHC8mNaHz1bI9HnNG1bJZqlhTqG/E7C/41Kwk/8SOxVvQdrqbv0
pod2g73FFon1c1gxOuvqNUMWZssbRQ9kEzuJXnaAyQOnPgwG4kYIo4ZtakdFtJA75a63QfqJVnB+
HY/+w/X3j5UcW5H8Q6f/A/STJ5FNkUevS3CZurZtvMim7yO5FNl26BZkudbjzM8CfvasACau57kp
7kgFkDIZw4u4pE+3yuHmeZ4TAThoyUqCm6SghVTsVmM3Me+ACPVpRgZPDetmhsLNwDtXc1wepYmj
BgMywbv0fdEvSerA5QBI28dJ7TyHQOyEtC8w4DWjorh7+iq/uqgx0EDJs26lluEDm8OyBHrfoNPd
coly127pxs55Nik3QizsEFcXTHLAKs6a0i0xAUE5Ybz8xRb/f5OqA94W6VeNqQSmGRjHZ6obolcy
0KdJmYKFgudvEHNs6UfEHADl887afqyrWUd/mFwlYYovIERl/NFlUFgL4c1+Ii7Mxt7WTKREgim+
awSqOJiMmPu8TAz8Iz1tkpH9q6U8a5N/t89i+3YOG7R8XHwxS1H6Q8TEPOnngjXniHGacD1eSxnN
+huaWgrfEc/s4otECMo5zQLdcBTQS36/YWwnqClS/EH7crlCgNtEhXd4qdFM8YLXYzGQvk2cRJdX
fptQmVTyWUL70rRlAclJN+IVXMCyUPIyxGFUNpBASUNT2UvX6RtNMis82D3pR3zxyYe0I5wrJ8XC
2Yenzetfim67udX2EbxEvdNi6tfLHfh1zPy2e1REAmAM4Y8tPoopptAsIk7ZNrn7PyK7SerYdJt7
JHoZy5I89LjcMBBXKBOdCnJCVr1y7Hv07gQWbpBmDJHFGw0I/BWsC5b4uNtbxBXbD07vu/DbzUju
rQWJwCpGRVTXhuuV0wzUfe4lZXW4nNou2DA2AzjHP5E5Eflb2IYswh0Mq6T43eWa0ueUDq5/we+K
bTdecAJnVbFeJds2mSBCQ9HgezT7CVqZ2/UIVLZ6OSp913A/503pgI9tYBUKlvxQl5yeXgL1D3ax
tyMXNeU+H4UojhyEqFmnNh/z1/v3JXL2j1zUbz3ZTNM6cZxpDaSalmciPnpyfscxX7rpXqw2hvne
A7gPJEqyHMgOJJ74s6DVgl/GxuGQy4tAMTdxPYNy9GSfm9WNIEu38tpGRKFVq6slpwkrMuxhi2px
egDh7T+ZQ8u49LK1yVA7VNHmkxOQc0q0qil1Bh1OVsiJI68LAONSzKhxd64CW3kJjvkmnoBnuf0F
c9aF8T9OB7SwaaQIx6tPv75PNeTatBUoA/Z+AsNsC13aJQHHCkcFLqeCybvBPG7Zwin40enBGK5J
qujPnOQxza8UWmmHlG48R/ZibUocf/wVJu2SljmGuKTOT1Dd2Qik1/GX+tubgto5ipqyWR9B8BEA
QU5EIqJF5k/jzmDhxX2piogvvRHd26bJlQlTXcpvmacAPB/AmBurHqrkSE5FpAicU6Kt8fSk4KkC
edxtYFqinAK/C9cqog765dpQiEcuwjUUFNCCJ+1w/3kbLIJlHXMAjxA2/DOO/+ZV1Jzvx/PHvTnZ
vD7hA6GQwzc8JPLEpFYoFGQtXu+nQCHGGncuoiXAGD0d5Np3Y636S//jXCOsXoygKoic45fgKyOy
ZrFuDC/liAUhgIIfViA2PyVAZVpUaTtd+rAnDzLG5xWeO4aiLr9UPHU9KqwZ5FrBCwtROvRmfRNu
NyRK6FGVyVooto7kCUiDbziBQIkhOf3buhnfpIvZi9QzkKvXsW6mTa8d9EdEdZOeukBXz1KB6p0W
CsqcFApCiZ68ubJDyqAejKmqyqtZWhWH09DV3kAsxAr+t4bBELVlbmTW/TEUvi4F/U7DjenT68x+
7cl3VabNjWUSC1qU0q2OjGsMuFWcyg+VHLZKgaF/dei/8p9yGTN7tb1QOXvyodZD97Diu61oyu8N
6Z5sBXXr6IyNdKAkESlnbUIR6TweAc9VWhpSN7Qe/gOfFaBG8aLbmZ5d6zW6AqIlQApoy5jZpdsq
txE2KoQT+VhuAelQL+HDeQ5OOITuDIz+yFGOodT99zDp/QBmFTbUGo8VDZa7zPtiT+aOi0tqh4vY
SuNHOTNSKua6rLBmvcj3lgZf9Fw11FAYAHyuch+GohcLQDk5i//JPJ3c+66TOk4G4mSrHcGd9EtF
exueM/QZ5UAXznN8np10Re/o5td+viRo32CUAk5jGG2hf+E6E0ZA+QNYvhAS8NmB98shT6bSH+gk
xjz9nMf84LKe1zE21d7PXO/Ow//PwUc7gpmEQx4QUxXs1KQi2qUOmqd4DhsdQdg9l15NKqBh/KoK
9Q1zKbteNTonHyF5QuGDUMa26HbjOBxF1yAGk2jTqQNGRz84I4dqpTq8hk1rWOPhVhtl3fy/LKQU
MKOSEyIA+FYk9ZeBbc8lXCnEgNBUG9R4P+a5IEC6Sof23C3RiVrZxBmkDHTshBZMvVn/k03+H0o9
OyBRKXnVlgUZmw3zEFNRUlnWchI7jWGe6wnsyi8bNXO++xCd4ilr/ilgEmudxL+HXueGy/0yVQGo
Y22MRKYYtV5AH7HD026UBTpLFUJieVMgE4GWC0Nayz6rx2hZMzpl5pt4HqK3Do1hrOEu6Oea7Ls4
LOsu6hMPc1QQzB5CaTAGgoSeXJrKs1Bls3CKF8ZdZ+gdiDO4OfiTm6w//e1SRo2h2nvCwHbw3C6N
WawOSlH0hgu3XoLrbtAXofoUm1TUAo0iEu26pGsovipR8AcNmoAsC73pY6wUZVEPhDWLP9Im+ksU
YdTI33dk7VxkN+aG2+4uAI/YgW+0R9PhjQkyZlDp2dgSzNZ6f8X6zbjdXGoioYNDbjHDXCZqCiYC
QdoTm53ymLcTTpf6XBQLWSRoNn7OzhZQgSsde5QBBwfVHlh5EgU79b4hgSrACA8NzCIebVktlv8Z
ax6H4EqECWRgZxy0goE9cPPTpiBCsxbEnJNRnfUE6NsHfJtur11cUxYp8p1sPpv5Ef0j9ZJsoBEv
pEw0yY75cfv8UAa3W+iBAF2BDKGcUi+5l8jHQvLjo3qVtMoU0sL0JDpqWSaFDqEE8+thebGK+Yz0
mktJfT2paZZ92TEQZyraE/bzx09d2OanrMu39kXzkk1o3TF+31F5dw383sE5GeohcmTBPHmU2xOF
rzG7X9L31SKqDKS2+3g0PBh4k1iYnrEex4OhomO2W3TcWr2qZe/EjKiWSvmdaYLp2i7qlZZ9TYIK
K4zEPRdguvAYDmVKkuiOrl1vDOrQUVyTFGw4gIHgNV5YvCItuP+Kz1Q2qsucwODA5j9/L7bYwcdI
awuihbAAssDBVNDJAmSGwff/Rb2vKHI8ltXLGNaSFnB+R23xwrTGi/JgWfs7vFdxVeXnU4kDGQ5s
uW0pAX55w/P0D3hslAHc9/+x1ciF9aV+saKPBx1Lc2r26oVR8m5OuNEwiFpJX7pdzbGs7oIZBYTy
fQFx+6lD64pLaqly10dUPFXwcslzvawtqaOjUl0YiX0bJ5+8ysWZHeRDby33XFuAttvdbEZ9HTFs
uYDh+WvmR2JNgc5fwPxGb8drB9Q8ST7geB9GRlcFPt9PTmeD3iYaLCTntPe2hCE8ImW3ggr/VywX
o8eE/R8p4tcDMvxRSCX9qBEetOsR16ywJwGsxUnHHPebCUIJuwBVM8jR11rf54PSYVJpAb9Kn75E
XI+JKWd1b1TqMOb+M2Px6LTFJ44DFBvcU96kUEbbX4nMotuuKTvKij77v/rWqV7c2qvb9geQCrge
ZH/ght78112J+4qmc2dU5So01Tr7MEUINP0CHPuYg99r7RCBMK/KbA5c9eoOtLvufhtNSJJJXzH0
CVpmo618BODL/0TB6Es/nBi0beb5kHsx2IFtaQ2Q1VDJ0CLWUKKFdcneSs4pZBVSJn8CGAi36K0b
oErO6kTfeyoybcJBpJ88EFoRzI/ajx4hxZbJQpc2AzANnHjHomTRsmIwNo37rE1ux5brlpFvy+Fz
4AzHNssti7N+bj6ylHEUpkLXEHD0b8AAknQxBuRCz0U7IWlyt/GmiETPq835qx44ZBPOnz27RDit
cRuJpF/2LEcGBa7el/s60JvHITSID57FwqoDk1jnzOAkm352LtEcXOHF4ilLrG5cFf0/+7nRXWVJ
z62Ce0ckT+V/IyO+GZP7/LMRcYE8iOHuZkKqJt13Vs+Or0nyyOpLFgAvxyM17LdSX+1LmQoXj7Ia
fSJd2dU3elKUeJ4KoI/H/k0TXLr9IZ6ex+UuH0mkFEXYFvAKV3lkSaPkr0jqYLzG+zWf5FrSjwVD
kvvo5P6RVV82CkVYaBzrkDnAP28Pc73+dZam5RfoX7uF5ANjdATIDEMUUn5p3kkaN80NO658i7Nk
cSuN5rJMs9CEOxThhxd+7ren0ume5YPpPxB9qk13hRPDBIWr6bXNQiaOK8IFtPMqBM1Hayh8BMW7
5yO5agUe7BDAvdFXP6HR1cshhB5hlGcMWnSOSpTRpbwvB/oiSqBCjexfpOl/UtifHANM+8fgyv9I
BMrX/LcUcB5eyCT6SSdKbMotz3kyJsXSp2MdysZybWZp09LN+HlOaFlM55Zbb2Ve5ELAXDhxIi4F
WMf8R+DEzCPMkTZdqeB8M3AByDu0RO2FvnHSnu8vO8ro+6Z2jdQD1suoJ6epk+aTM7NGXGK6ZM9X
XUhUeAO3y5/I/bidf7k12ErJsEsbjsuY9WwNczgnhNvJIpX3dZbKfnJils42g1vm55+dgWu9eYUc
BBBGFtm2vf176Ndsz33uBSCnhRpVe+gecz9Z4J1+faMyNZR93LBhIgpAL7mZDPUfMFLBUpiTGYkG
zkyFe9aOGH/IzmzBMcvjLBhjJI5C1xMlcJitD423lzd7BbGoKFdRrLr4q9X+WP5HXuYWycUNsGyN
KXgNmFuFaX3A354obNlqIZxP9tBF19wWFizTF0m82rHQXMGY2bEybBoNG0KqsbP/oUuaiQrKkzRp
dUDL4fd3y2TrL2F23xWUfrY4pmPxrum2QvOZl+UVU5FZC8ou6ETLSFmfFKuTGnWEKS/3MppWdwb2
ml4kd79BPGs9NhQ6VwgAgDqdgzfz4XYWeUyVTigVeJPxf0Oykr2CQhCH+sCvspzgpQgdQPLl/8XX
bk8o2z2sKi415nVa1nGfi+8gsGQpzFqduh8WmVjypQo0uQV/cb1ntJIbNtLM4L2QhtLfUQAjcmRe
JhXTx0GeO58qGt1nV68h6T69yxcUn4ehSPMdJH1JzmpPd0bnnrkJDGQ7XwVzonbwecxy3r0r2hht
+B7yEa3DyTbjN9+vf++u4xIYuR0P8V9qAj0IzYQxtIKuHHcqgH0+QmOPPhZ/yG1X+cP8Ls4LA3VY
zDp+W2MNjZwKn1nwBFXEdP8YPzYzD6+1i1Z6AcVdHrZFgnFMWzCHjLSxakFfuufrzKpXKmetW8w5
Iyl3Qumy82ATIlLX+bxvkvXfVnonPWwjHtXzD1EjW41Ll46532KQU90t2BPhTTllipN76rnF52x/
JnEu2a2P+uboX9wrzBxxQ5jXVX20KsfvQ6bXkIumj1iZaoTSwVLq15KcsydrRpIQSnAYX94MWEtD
o9OlTvVOWdSzVZKyYp0yMZ2vp/t1Lc7O6/UV7x9w/USNmqEQ0uPBdJf9I2DUDcrWD7QQu7gnyQlm
6uHtxXf1FoDL8183BeXLqfzAtLGb7rDgDPHj64e/KX+oNhJI+7PneAeguLVIvtRqnoY45WVRYZoo
7yOyutArG7bswl7aI6YptSUv9C4VfbRykVd3z9xfg17iHOtJLSdfQ4zE9ukovLuEB9JtXdtqP6jK
1f2rz3xw+yLGgl95CpYDxMpuFa8xICK1tTQk23evqgzkYREGZgReAhg2qKaKryXgj8gVCdqaqpjS
Be83nrr8Mzm8rdFBfAMF7qjXaIixKdeOQFOkOeD5RRq98asq4oqvyCFaE7+bn7vOqjof3XrPBPdN
Wqgc1e0x/bo0gdJr0y1RQvPiZ0C4d4uVrl8/nqBoWFPXFtPjj2KhNpmhIqFa7loW+EmOx0nsCNul
ewGneCW/gElfv46liU57+2ZX4xE4xbC/615xldcjzkbn+UnGMVVWoCfWcdqnoej+eGGeYXmdG7vC
Uc2AoTWNxdk1/s6+0QnN9kEmwVN3WB6tiLGuLDx+sB+wKjWrRmA1XTUw4KaUpNGrTtLNH34Ep+2r
5N2vYK/g5k+Sb8aW6+p1r/TanlhJ3ZH2MeBu/tdZTnpeixa7mHbgecixQmeZpYCyQ4ABcGeGRhII
yoyvVYeKCOZawUwGuDxDMY/ZbAQ4kfkSb5T943XauzFlJjSVXm+9XP2m6cp+Tde7zUw58rxti5w/
yrEsxQNh76Ghg7DguzmomP1qMwrQbguhZhsGne8eqeTN33a+QBIk7PeTnkdUdXgcyaZxaLg5CpAR
o0esnvtivyQkAcGaE7xHhBrUfisSCT1zn1MB1EGvNR9FtRvGrEdl3/EsUyIJN9cwA0tSYpCBdgdg
qDTnWRSnSma8gTtgkKGzOVIXxTGF1MIvt6fOH9r+bmyvdpNB+W9fcsJYz5TVbo6AXeh67Vp6Msr5
OfYdDNVe4llgbPM/HiAPaV/CQWDTynJbeYWv0l6oUntMRwSlg3jvQwvqOr2n5pXU56Fld8qFMTtj
i6CO0MbeQJFTws+vXJ+UZMVR5Vwxv1t7LNaF2bL++Mq6Qx5oi7x6fVg6v0eakXDI8rHWey+fD5Rn
E6ATQGlx5ChPFJTKrAAbrGPimX4mVnJ8/s48ZhZuU7vyXXiDxbpcfBkkRMYhHI3PD+tFjDv/VhQW
x3CCfGVy8ecWKSgqIKbmFcs+TMSzmvpacthbVyb7Bz/V7JebMyJQslicwMTms4sNielnFJrI1d2U
8bhA/XfMLSmpsLtYZxpOm0kJmnV4Zm+RlhWLydtxx4+kdOsBdcothVWBbvuCAADHp7IRpHDXqCuO
+r5QOLlKrNUDS/lu6+wSwPYINHEDzs9HDlJd97bZT4Q7Th3MAwi1RoZz47mb0A56OnrSqm0+cifn
gWP1kRF++xf8IGvIq0ukUrj09bUhcr3Oq6AjgPuVUXuBJ5j/6zR2w/C4ZxuDdRRfNDKJ1oeUTLjY
eHD6zR1jQRbGLG3zMHFf/7diBK6jSyIFyfwDupxwC0J4xHXNiu3Fzlbs63H+KlMNHENrftH+P9DB
qzdSr+ibRjaLMoxkkrXT3DF+S7uVnjdMbqqz19ooNJNTMplYj3DqggyMV8dKhjDwFXq74IKNC8IP
yZqqb1i54o5/A1vnBJiD22arMz9+UUqPDXPT74MRYRfbXppnL6gC5MgMi8MmiGwMQ60b/tsZbDCO
q6q8niV3VgAB8B09jXd+myevgS1UQ10wgBMXwZg6yBmfoXaSYGOHgThlhLBepB74gsAvWQJqwxR7
NDKclKyWgrB+3M/jz9xL/N4N+spdYH2JQXZwO8e1Piv3VmC5O9FvJhtvFkNxHdE+AyGQrgUy6iWU
CRkW5Na+uA1HF6WKEuS/ZDbczL5/SPrSju5ty6NpuVPSF3YtDR/9dG7QJsBmWFGPXwpw5dZal5+7
I3KzgzpgbC0wVlVbJyHFZ+hlwVQ+AHwgAuxvCfIEHZ52ohQtTwChyqk6BhQSCotGEEbT20DHZAXy
SUF3o4v9/lRBzt9Qku4IxVFLx6301MFkYxtTPoMQ3Hpzs07NYopH0t26bxG3xCrChHnqnOSf2arO
uY2LKB9Iova3XhvWp1QwIMDu+TlkENJRaZTi6xs/JEH6sQw/YeG+Pd1U0+uywjek9bYkVbDOnBE+
4DZw7JDjDCsB3VTfAMl86Y64NhwqSRdeOqWTHOlKLcfUDyDe2HjMVeZjVrWgLW+JeNIs330RtkOX
lp27AG+44GJOiTa3FkQAYJKuA7nY6QXffRlB6b4vKlm9SjRbjstIa/FXBm61cQ3ofTAe7SETiSyD
+zfzsLoGb+oZqj90cSpybZ91/nR7K56RIl/rnZVv8ky3Hn/qRKBAg6ck4HYDiySKIvrdIUSTXuVp
ILX9pJTXJmVsWAWzQ0wB5sZQjOP2y4Zdl4Yl1Me7XuWTv93CateyzYvRZt4i71ZxtYE+5teaAUKQ
T6MhNiaOO6ITIl/afnbbC1bxE9apBZ2Ha+9B/mRjD8JFdnpDnidWqG1HyPeYLQ16R/TtcREW6xGZ
sp8Kjtp5Zl2JuU4W49S1RXv/jzikEp+Di/up85mZ+RLCNf+G1myDebH7aaew+lqef3rUzfBCQPjP
r/2MPegzr8sT4XzPPE0btjMfEMExF0XKF405EkZh4aupYAmSi/a506jcU/leo7AWNevJ64u7cdre
3xoMZQtuLIf9iYseABhbDHBhA+jixHzA3TvLaE3FxA9bN3sXb4OVYvyErutQE2m9omxzhMQpx9Ip
b154cJecy2OAuF6H+nSqFAhQO7qY3luCQhGt3qnoiF61j7W5ejiWj7J12OcvOKmfArVGAb5n8fUe
L4g4YHiqUt8HPPOqy3Q3hkpGWdTMex7xs8peG11kI/dv/i1rA5f2hXJrt2TMSOhlHhlsti6OaHIS
LPtRBgiKRIjtOuYUhhgOn2Pem9qgeuqYum4UNfhsnW7gAYWHdmGOwHfjpvTFXso8+u8dYmAF34s0
wnQi6FFp/QVw1fHHkdM+77nq94XNI9tuBShCVrz/np3CcdKbO6HG5PmRtzBsZxDSoJoI0jhY63Pp
jEaQ6h1psyP3APbJypWKQy9zvE27namteQLE9f3KkC+ooMSi/TYfnuyaRCeThA3k1Uu7FaSoygUI
bq+PgneYLIBkOL+Ux1BFigqZqAjwx+nK8brAhQU0A64REBb2UpN5nyFiLRul6A7EFPMmb/9OBd5a
xL4yeSMY2qWS7zJ5InjHuW21shjJABsus06qHYyH5SbhI+STilOaJ5dRfDc2KALd7mV8HJ7/lH3M
NxeGTq/m3Wr6KfsKc0+H9YKEVVL/xWjLif7419IoVBZJeLJ0Br6WbsjAJFDtM4tHoMkB+Ya/l9fc
tlW6H60SqvUkKiS+aoSKOok63+LqsNndXdSfjr4BTpbTG8QDz4lB6Spz72u3NhGlBhVvVUCUQLah
4NNhYTD7KCRmfuNlDwJN2mioG9K/rzceaQeUEN3ta8U8bKJh7OA8SFUk1lrJKsrJgnTtODG0U0fN
ZRkn4wzP+Hf1zGwThZqIKxOd6NMG4d0rndMcjfwVcNt/zGqynCmQ+oFyFbe+ujZG2QJFwqopAPse
JTrsZmKVxK/k+SErBPu1p+2c9KPhQZiM8WvRkoJH2ocefwT+9wGDXSVXf03na4Hc33BXuDLwwB34
pH5Dr4xorTWbpF6oJ8qNyyA1SPZv1O+40Wix6NXRePtEyFe/EEE0N64RPvtrtQrReyfqwAx7P86r
uIaIir8PsFlgn7Oqnq9+ynUTQfdjvJO7geWO3dMKoPYf+8kEOYwy87Pe63tVyfl2/1FAkObea4Cl
oAUa7WKgMblGRQqiU4JlW2LNXLiURZpuvahfTP097mC/qhfbB8CzellSsmI8fiWDvGK1uryygRav
GiQb1IbtXGOHAxmJQLiCzPGrsb6XHRHSYU+6gz4oOsZ6mMABdZNVNdvYnnn0xN0w7RoZzCcMPti3
qp24RTARN339zMxNx/YlQ9jESx4Khr0XC4JqVdoocTaThwy0Lq5t7AhSZLdVpwpEUHmcRynu/7M4
I5cRQXehDb5lZqNmhLHZST9acZtznAk9aplRRUpqQuY4Q/nliEmYrES0ZhwzEb4zoTSu+cASce6s
3Ks0nOR0/cbLznwN2z40lqrKECvmBKY8/gbooUWTyYzC+yfyTEPM9A/cBEk6sd1PLNkVT1Dd3NDM
LiO537aeQvycVajQvOS0UmCp3K+6QvGvSV7HttZlZIgVmrGhj/RXt/hue2HLKfX2nJdt0NVtfih5
jBWntBfcog/c3mAaYGYzO1vZ4oAXcyV2nmqxx4DpLacY3cv402vGEuxDbRSCwvFsXjWZake85Hlh
RMqD62Rd0Nc/32ZyTdsnLZp8ihaXO9SZkx8YMySiY1yCuAWKBDxZIirKYgmlweUEsSim0h0baNuI
WZpmf1ZPgoeko3dhXj7WOFgtgNtd7tnVFR5sfzbM14TXvlJIB0FO4YX64YJZf0elocbjFlEBPJ79
Cq4Ggl36hq8xshzTZOjJ3NX4qo/04bo9KcgPzWt0LBJCvxNVuWWZh/JIQbtarT6Pzv8OyKa20RXG
UEaIy5QSIT7fUd7bjfeWMmmxt9olaZWGsXY8HgONpfcDVSOp6zDV+1Ap2eavUsPsaJ5B0fhKymKZ
zYoXXZOszxk6kQBVczXrSHjQcLsuyhcvOmLThPRtMSqC/PkXpHuJ3AAYP2SmLykFxABfVRtDPgpQ
UuBlwKglFMEoxyp6sdADES+3M7bLtRuE82k7Yw43RsAHszmoNKy+iJ808b+1/4EixncjoMke2PxP
KOgvLcDrJV8K2rmtf2UfoLU0oc9pqZnpn/Dqg/IUywJ7pvif7qpbrTJARE0OBDvhbPCJDZ1sm1UD
vjPEUBA298OZRrALN1hOS+pnzTH8sZg5UoujW85ws8nlYJA4FPDS8Q3AGYjKUB1K04N/Sddx7e22
pJtj2LvZfz0WubqQCC0qSauWcES8dcVN072rWliXAlN/ExxcKYOqln/TQPuhEwbaMMdvYbJKzP8U
HQG+ueL0DSJqXkfJCLNvI2E56QHXVGmDNYneDZVRUheYj1OK/liguPnssUSsBg52oDeeBjucqHdA
N+zpDYi49ZpgU/czhTxDZT7hgmJTiMIbXehVthqiRJ2k/6Rg1NaGRdeOErGYryUlLw9urSAyyxZy
q+3lr9T0PipWVZy4ZJT7wfz1ySUK0a0LhXBH78VLunSKPwriZk27oMz8ho8wVyytiYk7Tzy+/PF9
9Y15WjtuFBjF0nUrBpjhDTNy7+XaDIKhhmx++lFtpxDXHNn4Y0aZOCJbZm48jS4l8ymlrfQsXTJd
q3aTznZuOXD1L644Ddz74fN4BPn6uItaU8mTLKZRe70E51BmM0JeeokuanYrLuyZeoIi9brmFN52
YjxozpH4J0I4ux52vOMpok9KdpApIayrPKKP3+c+2VBELAK1DSRIidZroTTzztXZD+WR/TzYALbo
Mmt5N9Vyo1EMVC9fbscusvgI/+GSyMx1mhR4PENSDNazndIteUCTh9xnjkvC2+UdIfANaShvQcu4
LXw/UoxdTCNikOwSWFw80z1O/akxFVFuBgnK2+TGfIoLHAeXmn7r0SQkFvl1APkw0oSysJyDKDXe
LneUoVh0OKNr2EXNg4bVAGsg+iPEm+PCH8x9d6w307qIFp2rZ/KX7e+BVTfrBPorqZdgpvHevlY3
NsCiDOcUcwocF6uK0vbrU1OYLg8VWD/b/R0n/ovIriou6xQfwFfXojj6teDJTgTX9TuF5opb+9O2
Qyb9FEI18NVmzV2l2tv7heLQxakja5zalj+/DyxIeb2idkkw5hzJ4W4mxm4/5PLy2YQVHD3W2oP+
Per0oVPntZkEHV5rm/fPHANZzhsFJgGgPpnttwArxBrfwjwtdUTK270rM1Hhbo6zMA1rOXF4r5J8
vI0QJ8RUFg8erYtviTZmIR/baRjd2E1KTUtL7BpXUnBONEzvx9PZqckvnIqBvCa6/y+dyGugJxWj
mw+2uUnOV3SwXja4qCTEE1oktfts6d07FMdWQ1ROZ3dSLz754I5LL8MwP0x4tHiDcwKqph66Zowt
bTKSmIsSvlH8tWJwAbSM7uN7vs0PFjZxzY4ygePQdktC17Amd9oABtj0N8jUnR2EE7yzbdb1XTKx
aajAi8UOUFwOJv2z+KIhy232GYr8fEvwVTKh4caJJ4DQzYlmRRjKRcspZNZip6cA4eJS7J5YaSSS
LUP7u68z7O0r8hnQOy5clIMjVigpN/VKcZvbyLqDcMCW9XFG2DhxRqs1vr0Jcg4Iip+vyd0oAxxp
fkCPWz7dL2WXSLesYZCrDHPBvsyfuuNWrvXYGoEmD2Lj3qmGNL9OP7/CoXyVmORbdHPabkb1pAoL
AMN/9w6rG02IGWh/Ftr5292h0yyYxNeo0A9pmH4h6H/UjKI6m6HPk4Fkj4+tKw04NQ6KSuX7FWaZ
/nQ0KQn+rz+k6Z+JTinfmCHf97rN13s/Dxa7Sm+yOGSuGrmBDoqDA4N2wYUa5G2955UNGybD4TjC
SNpMbLTC19knzwens24rQlIaECuA2e9RPaZeMruh6KAhn4XjEPhL/YefR9l8k5CIvhsCVn+Tm6Ng
3S0IjLgOBlKlzmU0vrV+xLmEQVGbRP9tq/U0mZoYv09WDML5GkSujFgYBJRgfd/lTs0fLxxFG/EC
MN/AYluEl9BBWnXZfPxNUpYL7FZ+zIfvBy+ZBpu6NHZOm55QTRWWqHUFQwq+nvkCFr/tCJ8rj66t
prH8K946e743wA8tQUSeluvhJVOu4Quh9UlP/zvAJatALmqOf0xwNjTlkp/DDL/8EKiDUHY7TVg/
Wz/PNdRQVd+q94Bed1zeX3e9UdrhqLbV+orVdLyh5WNcxZXAUauF1n99ecCQJw0Zf0kTut5I0B/f
McZkPe8BiyzTCloicmFRvunEswWrXe+g7zTkdN03oBGDPj5lXx1tX0qrh2eKh/XE7Kcdbn6XGp43
2iw1uMLgjqRn23wcgs/1YSLQUfQaBp+YQMShxvXHPSbpWuGLkPddJinAEspvXYBbtTKHm7FmPG5N
Ea4OnLEBSLWbEldBIvigxotLRpw3GrWeqJBqfT6ohLPl1Y1Q3xUizmEF8LygcMIkblhk8lQAdi/k
K7KJ/pWLISAsXetI6BelRt4chOY4S7PlbUdSltxRj8RNofVzZQ10RkpegNQZsJ82sfwW/DwkPq6U
4EJ8dtXWHv/g9s80zy87ASL/ELFplQYIAJu48ZTpZF6TTkUdJ0DzK2wa2s/uqF5Zr8D1/S1+CZoW
cn+3I8CEl0bMYCIF4S26/pMvbe9xC21Zw4oarAsV5P6Vv3bkI1MK1EBP6lcWxrZgoN31ZE6cyweV
Ox4aXT67FJJje4VoEvsMwgeGbV8kbtw3B12Qcaet1R2Ngd1neD6EBWEtHjTJ6WAg1R7JaPS3nJA1
2o0iaIE8+KNcAtNfTvGEHgEW7XHXvzArx0XmW/J/E1ISkvZmEVThTEqWfqoUV+xmWFK4Duoeqmp1
jQIfp0jUItiu6gAYdm0QryiyKszyQEBlYALcJXltFqeX0HQMmTEgVpNGo8Oo49osyO+XO9OsYox5
IpQKyNN5vSWn36Vin1wQCkPp7uokCITCAWrHKDj3KBsCB9qOSKUKqWGEPRT0x96xO8OPsPzLFM8m
2yFEwVt0RB4PQ8urKBcn9Noooa+MGU5gBuhKjaygogc+LhqSE/iKYbgnwGyc8O0q5fFWmhXN/cbr
rBCsyBPDYUwX2i43Sb+KCYwvbTUXVrcy0jjAQ9zTqMj94EVAYGvOZAMJcn/4dC3K9JFFDIlruDwV
bfW3Egjb5CocCr42eq/Omy9tb6JSgYHfXgTOaiY64JFAI+qmm7nCWt9kGuD7qTUlvTCCMr29lKWj
btFS4K6k6kOIl/VNKcZy0hESi7Tbw2IlGZv2yruS1jV9jUlXWfDFBQp7u+I6j6CoKnwhI0bfqohU
1XG9zHn0bPLtrrO3svqfgpK8coDhyD4Lq9lu1pAd+WLNBitmymf6t5Q9L1dilpunVvjSYKwQ15Mu
rJEL1D/1EmfaX4NZRBdH4EaWkow0CoTdTfp1V4KqxwbGGlQSLoTdIWoUYxsTX70RHrVttq5KENu+
m2dGOOY299FAH3R3XFrrHFktM8RrHNmt2xiIQNg+/0nvpDTs6R8IUUmPPZ0WZUai5L+3zMdJQ/Uj
cxQV9Vh6oxbLAQ59ZSzPzR0H+/TdUARL7jxj0YA1D3yeoH+74Fo7ssfMcCOhcCvUkjTeSJqRMxWC
F3vtZTF0leiFWRSwRsawVUw2vX8I+VErvfM120fkug8wOJzJRf1MDmDxLbJQs2fofP+EAFMuAQy7
PXO9a/p1TqpecHQR7Obh+I0si+MWSE4pC3GHiWLl58X1hSJYZWTEZ8YP4bXgVJf3GeU1Nj74wCKq
LRVvSWH9zPZ9u4r6nSFZdSbeIyB5blG0HM7n8DhgFEFcxSBcSaxVdT/A27blPGn72htYzZvbYYkS
CtMNPbWIuqHPqHZ0T5FixEMW4C6KeJKAMzwLxDFGHlcdA5FDjNQEbEcg1ukRAiGwWKyuT01QtG60
P51XIFQ5R0bEiQ9bm9Imz7rAheaqCKWMSN6SuDsxB+3UNImAoEoc5fk//CktPSbQigi1/ZAhBvlQ
lplnJuAqiiOE5o8UfWHd62Ov9FUJh5l8GOeYaPx8N6SPY4FDXKjhNn1HeuyBNq2R4L3WxNRjYG2k
r5UlKVMr2/4SDspA+uzQnkjP0JNEZpTZHBz1/179/PwNi9GwmnMzJ93C4MjopZSv45/bCZQBBFUS
WaPCCJrWGx7y5zoc2/HCa6DSwcBwohipgz7ig/+EwDkpXhtRej8YtlIpV/yFqQ3KGJuIQusz/qqj
LWUBNnyhQqjowFsRZ4+Wfk0kOR8pK5kku9QfaWJD4L+tu0nM3qGVto8ddG29p/kwaN3YMyvc+U/b
PFi14JjCe729/bvJ2sfcuAPnvMBEH+uXno9eyZTusTSim0MEpworaZmC1/2zRCl2Rpn9Lx6Jg4ET
jc3Avw7krKdB8MJPja3tYshVq2TII5GueyHj5Bd56N2PC7y8Cj6I0QJmwR+d4V1vHFdOeSFAbLMi
v2xu3bRZRZKTnHtXkZo/r6TQTyOMooAz5/+lTSt3wgcYua9k7Q91lg4Id029yfRBusdUM/AAPODx
Jkuv2TXXWoNSaSTdU+nQL5x1AsXrIuPWiB17wpVeUeKmRMDBBG44PqD5vU6rDxYePra5m9uKrEMP
E1BS88KtJny/2Sm88wNHMIIDRwvshB6GEkICjV4afH02016CZNtrXdobgEMvok9fTJH1H0c2kie1
8qE514GmIW7qWnRsAvjYql54fFfulq3fkrROMNNn7RQD5iZbLz634h8el03B2K/Vis5EP2E7mlQa
2QRycIAydhvt9wKqn82LMXkU8HfNiRBzkxXjNl+O/FJGydUl2bDyRrFJ7bnan/wjs6kx2QXalIEB
v4HRrLgUggYjOqJM22wdzznk2pNImF1BlEuLmjDhlnHTnpNaxP/jjzGZa68MyK1lVNyOBNTvOOPa
i3eW1VNIl+n4LuFqzlMh1SiCGSPWkl0WxXE6K+Jh90Flv3z0xcHCTt6aaQmp36wr+EIu2WlDaM91
z3KrCkghTrkj1hdbdeEsB7wxwtrXcfiXeGPoTILXg4ChPwXkmYsSaAJhvwCM1eXWtQjJyd5Kifvi
TnbX8krWx+fz5hygrFwNBd7mjy+Uu/QbZAXdRQrhct1VW1NXO1cMgTRSpG2TfZyAOquiswuwzNjo
Y4/+cta3L4Oxo+LNhwGsOLkatbgeww1l6go8ayoFzSsewtTzyPk7SROKox10L2DHeXF6UGd5ukCT
XEr4pyuWqM0MBk7HtSc8iBkVhRHhfX24qtA3Pby9kaxWcywjgFuMoam6Z7yK4s6kTFf8RF6OnF/v
r1D+Jh21WW5kDqt0dCRuqEhHqGg2+N2nry1nmX0lrYIAOjpiIoVV8YxIwoC02Uw4KC+GA503jt/N
vMMkxZoj/PypnmymsKG4QvVbqntKd4vwfNtlPpSuUGEPxY0LhZYPlXBfUL1yDgHUPwEPFN4rFKFy
vz/JMO5eDo0njUXpcn+5Zx8045PM+m8WHqf8INpzCcVGW7WXpJgODKzRYLXfHdlSgwfiX8sYaag1
dD8jzXM511F2tLZsJOniARMPYIv4LEmzF6qGjRlcHQpk9eL85zeX8uQY+pmNYHYDBa6Jqbsxb47A
XuDeWsUsqNIS4VkSDK22ghAxIpKhiLT9KmuN+masn1RO4/NF4lMs8h5XGbkuf4KfIdMY0wgvWSzg
wtfg5ZL/CZmqGKZhIUqP2AYviim5gTr20CHjDJ1lU0coqxshnoOtVHI0O4hwPIkJwkxUl72Ku1aQ
NAUknV7TFrlTGEyNWHkD2DYukp7aoN0I/9H3/S5wqW97GhHOl+sBLQvClYrTtFBh+nfIs+vyAQNt
pTa499HNY3lII9TrnFHKxTuBTJh0h60jGcv/yhVdEK6CVzNaI+AgJPn9KwF2aCykKAbb4l5SetEx
QFDcZu2nOLVTl8I/9aVobC2gIwGeovMWHthQefJDAVT/oe6eEZyhZOQ6M71Uv3yp7s2Fmnd+2kcK
8m+c02V0mMls2M1IVwUdNwKKUzxw5Auer7RTKXjRZ7RCY+13IievdCXgHl5bpJP/VlHPqMwGQsCF
6pn+kSJoGOer93LyxCPwzGTU3Xyn8fSDMskhuFyj3y0ly0u7DoByEhjMSg04JSMsmqGupaWufM4X
sv1XWp2SL2t/QoV+IEt2nsGR847Gz9MCl3B28qqkyZ8UykTnHktrSp4rFNbGHHGig7hu0SDSASTZ
Mca3yeyzAXI87e0W8BLGTIpkGKKyTySaogjtmE3msPrKE+66jzuzAMOwlxieTpgLCAwNdLqxafys
t/DkzlS+tver4i4b8T3uuKPZLYeTJe/toLZ1c6vb7QCWZxEEMi6cH6B5Ha28Exwm3ZWH/9T8JDnU
I5y8GTflhzj/YAorp8IZ2Tw0nLM6iQHvXd4yO0wgwNq49kV3x25lyPLmj+DdqHiuKML2iE0OzYlM
MVn4ZzWLDMhkyi5woEXVfH7FKzCvcKLJPeTZsBMOuXWFPjRehH/q5jZlchnE1WFNPBVQL23A7G1Y
HzLSKljI7EWpptgUfqieiasb0X597RbmGawqHf1itktRx5eKWaOSotUQnyWgPydSyIfXuH3YsvIn
r32BbH1HpnKdeAs8dA8ht2wp0IOPTJcFXFB02xGd3g2/jYR5rSm+C9+668G1EdH3k907NHROyUU3
jvTeY6ghZwnmsi7C3guZ6r2Co8t/u+WxequNIV30XSebDF2i5NMifRMd2ceIkaldywVGGU+UBKks
5YGaPe1dXpq4rygIiulJ2o+EoZCfkIiz//11TT/MZEBY4/7KF776O34DLaeihOq7ngfxUCCTwCWQ
LEaa3Jh7lA/qUhISNKFYCuhNxduRG04gPca0gf9pAmv6c/roHIEEgiYa1SMbOKsd2Dhu7aeO04rb
c7Lcp7JGqxXTzr1h9/kcBqAEb03nFoufT4dBHGtPlwc364adRC8okzkPWQXAGZHHqEs8GR3Exzws
qi4PiZtHGB9obTKRKFYBY2V3oYkwEomaIMSCE/E4duj6Ms/0QsTsGio5RYKyF1rcM9xD8B6yjGbF
+JtO0euS1D3yGoxgvCsA4kivh6/yinweI0NXROAz+II0/JNbQUcznq4tyrUuDOaDC4oDpUd86Q3W
cf1lEuVSgyCuFLyYzt31fghRTLrQjszu/3doYzHGZ96iYEcNO4VqjBIqm4PLLnAODJ5ILo9QFDju
0GrbtinQQ60UH1EQHUXuTGoDEpn9Y5UjOg55FkS9xZ2bO17sQ98si5G+81WiKKx5By/lnpf6r6NA
ywDyvZmXPF47iMNLm5Z3sHhn+2pfmx1WYDFlk2XdrEi7V2wSxfoT6MMDr7M27EpIE02qLcVV043v
bsMj3ytfeAXUzQstRS1o8lpOpTuQ3i1Eds54JQtVqWHP3EGu2HbIhiZROF2fB3nuguzr1VnGFfG7
/UoeTg78DtQjFjJY7wQuq/9mLBw+G4CLr8/mvl3xdHP6qiDch2O/trm6NLFdEp0Quieapd1EjNHR
/eCQfM4JTXB6zkUUiNFao1/PR3F/7An7fyWofGU/G49WB+0durb9UY7KuoVPNahi8yKi4PrAFO4i
kqlIVtu1djy77dnfoBf07UQBgBtYFqIb9H7IahKuUIYnox1pVP5BkiKk10zHr30VZAQCVEb4vEFv
YLivYgjDyUhdyjhfI8Dl0eC7oK6n/DD/5o/PT4i70njfY8eJKLYCMjGV+VQthwofjO2BoA2tlH0q
+nEekv6PC01998B3zDagD55tEj5w4NGNHvAwqD/prCt5/JVIJoNW9MFHopYZPICt8ftCNXUBQjzW
PiCKEv3gs5tVMq5SagujZN0z7qGJruA9x4Hn2a6vXKCs30dAHZPyZfsvzEFxW76l4950NPJUtRIX
0+aFl2hwa0NvSGZn3/bobB9m7oy5/+U1Ar235HLJqS51MLy0640CbefqTsHfRVwTuCT6mXf7A3vm
pKzENCeJsdpiLy6OqJfZre6w6f1z2z9qFy0Klbx4ynJ9bxxzEg2qfFpIDElmu3xNC5a4VUelzL3b
m5ubXGPKhSziR4TEp78KQKcsGkvJJCQL4JwCI2jOE7pRrkJUyShZA7HSqNdTlP/hV23VW5/Tz/RV
u9F9by+hz/Rsy5B9K/+Hk0H6uvKg+bfXDb/VYHW/dpUcTPjdEO/MmoCBdhgGAXxtTbg5Vc0yrDqm
B4Z1NhWM2UevtyY3L5sFAlAW/aVrTK0tfdq3j+cXlCyj8GnxZpypsBb+4/O1XEhpDjZt7JWuSCAn
qWz/0nmRBIrAVaYkVWXYv5bqRjEIG4HaUlLSFG5ibKbZUaCfWqr7sPWZmZRctFQAPPCwc5Ew8jrm
8NWgUElU3qL9DpSQ62gUA8rqZR1H20K2/pRScu/RlJ5VG/8t6rtJXzoOUrOV5LrH6+O+2aqN/A7W
zB39ueYbfjV6jdu2z29f2BStsgmGsDMgDZd7h2KiNl8TyMEh175SeTs3d0WJf1GY8JNsRebD/r/L
7cvfOxsQ6Q/ekNiPJh13Je3lxatWC2NNuIlsWJzVUr8Yvqa3nhw5bnWcUgvX0U2ZuX96axckyZbW
briWm7i9Oz6UFgEPM0KbHG9DiHFBrzeYVlIF1gBVBODDjWAjxxs62z6ImmDMwFSJk4GnCk82+iml
X+5gmpY1MQvFNSPEnG4cXX8kYQ1qNeulDZySSKwmZfU0OGj02hPuoqdCOm6hv52NGblPSieauyod
Z/woGZROKXNetSfvVX380+0q5KlKaa+KnSTIL2h8eKjwDI33lABA/VypzOlEJRSKTyJGeWtjQ4j5
YC9DPJIpfVhlGg/VwDH0r2/xhCvLieSTT3NjtnCcBMo5g/WvkpN2vgEJnmDxjxiB7SKY38xWFV8j
s/+bcFRWDxHzJTZVKrAMPhckLU+2TeERZChxv2lux7VXRC8FrkbBeJpss1uBcHx/Q36CrW/hwhhL
uz2n98P0Dcczp1lZuIEdgJm1YKK9RA8xeq5412M8umD6Lpay+X3b2rrc/uUcITcNf8Bd0/1xGNPw
Ofk8iu9q8glUxdcvZMnoYlLbZ0l3L8RGbQxu1bKleb8kh3l1GBODGmSh6QKechSmfn5g0gECi36j
NOD+czcnlRK7Im3Q6I8JGhDB8jpzGQQFOO3jdElW1RIdgrq8oThJbNBhwmv7itasrjDGJ176vptk
vvo+TN23MVoznhefTKBN4vNoLJi9H5XiXA51gc7ByISItg3oTu22LITLN5ceXd6FerJpu9nVqma1
vVYqBoHOtJmqHFswOEnPVH7weY3zv4lA0oGSvbS+CcQk1SveMIm/oXXg1fLgJ1DAVxXlIF15c/pd
44KTsYGe9DouZf+wz7b6x+VbdHQno+dFKEIz4r4xi0kB8guPQehovtPdfbstZrC4y/IwC3ZJvPmX
eOgwOOAKHU2UfrE6U+U3CDdFkvkFE6j3hg96hw4iY4G5W3tDqfzCXeOWwWaAhfvW9FprYZrxzwmJ
egujqcEzjP/u8p5OqtuoSQEZ2x83IgZwj9qFUkR8ZsMTDaFeDes++zp660wFjDXk/qcTXNycTXXA
UMF4wZpkgRxdTZW+Ip+UVXKAAt0qepZjE2TUZi28Hq4SkrSz2VaSUWEgsnZBA49BBMrANHF6ewDE
5BthlX/mlaBZBTW8A70psatkyTCqrU3rprwgpwNRiJvqkcrBEWKcTd3VMcz6nVcit8pPQG0ydsba
/djdodU/YIJPUyo0lfgqZkv/rqrcTu4bvWBD+qKjBqXkUI8dkBlwQNGTq5qnEMEMlnoTCUv+jK1a
Cv5LSVHUGix6kzatAtlPITDaEI5RkLkpXCxvlmBwsO0BPEzQY2shwJohHmBLqTgIEU0j0If9WHHY
HihDWreitwp9cOoI/JSUBfh+LU/aBuktp1WvqJwz8vtmK8X3FyF88hNXAiCrfGgtomxOMIrGjaFM
jmSO762LYtyBqJDLe5sxs8rkw/OXytD/hmXsthSa0NflAW2OA3sCxInfmUS69GipRNdCe/IQf/ZC
occtXAUsZB+p+kvCtARR9T9Aun16/HhI1aewKEx/VmY0GCOVI90ayC9SAjIktbD87bXhnRdl+YgJ
ZExzux1krbgbVrbNI2AwPzTMT6CRrDhqiJmdzcaXeTqPOTMUXcy7JRcwJA6rtTXkRxviefx4kl7k
JsRcn0g0tsEQoi8StbDdN/qHDm4Qk+9wC/Et3gYgz4HFAN5RVBtnEtppuoNZxx90FMRKYK5KdOpO
4TEAK66UNAH8nINHFGMit5qen3KnKIngvHVmcYnZP8Rg1vv5VBna2h7Pz2/TGZlmxlugH85iM5i8
PpG6dFDdCvkUIrcYgJc2B19iUMVsxweMZtOdjzPf0f6iR4khqPs6HMCjEit5uEWdH6Rokf05G6Nf
Fnn1r89iSNrP/X1HNBoX1IpdEsw7keqg93IyVXXIPGmaK5XiwH8oRaxD1NbsvRwdyN7gBxntL4qO
UesOmrptfru9yTZ6sNK/wgox0OkmXN8KGjiFIHzG9Wj5zJlf6eufnzaXC25WarLvgMwp0skBDVzH
fCwO3BzGkt+TZbPlJtirwJNuzhg1Lapq6sxvgvyU+X5rqiLssveeEyQgpvK+9DErvN/Or73Bwc/9
a0eGSJ69J/rBtqi2JqtHaPqMrOXQaR9kDVoYfDczMIVYB5suuyvBEiaSA5einszmFAIJjuu4OhdS
MTkLhcGRBRI6kux06VLMZaOtYs17tLwtlIfd9QA41uMm62mr2JHVu710eT5rteJ8rvuJQkq+x05t
lUI/eNRXgkeiRUZz7I1LEu9nMSKZV4SPFBXzgXXK/kw/iQuXpE2rZXbu36/4WH45XHKXyxENLgW7
yPvpYXpwAKtkbLVXORBzeeGcHFdKVEZDxDzV7AYdsqUT166wweaSbz30WPQ797x0iRAcXs7QZlZN
v4Zo9ZzhJ/AMxdaGZkIKTYK4rsBJQvOxw/35jycUeejZwCqyOvN6O09/pAZUddehly/tKC/D78qi
MhYu9UKUvgJUu4WD6cIO8/QlNiAR/jIQpBxOMHiFg2qgsFgmr5iDTd7sr4raJGwWu/DPmwfNDLvu
lvIfLmjMdVvTIkBCL6u3aCK+AQwRBa9UnqVPYlt4UWQ1gt/t5dYJrNMa/PwkyqWxHM9UT/vRy1nY
xDAA9qSwSR/4LgCRmZfy/XRxppQ7vTzLbxnXZ7n+HsVJzQ79y6KfCM3nwAJz3xxgYUvyoC2c7Bnl
crfXLLjmLRlDCRWBHjjCt3xV6M32DU9nfYtF/VfuSvsi4jl8ALH1oS8Cee+YBkEMPgkKre6MIQ4u
ORGkJMmTyafphFSbbxRQVD7aDVSXDYoAZgAeTVLqf82AxlXAhkKJ4bHAHFs8klWJIhr6xEP3QeGq
mgquqnaWcHc+hLc/rdUPZyRQ99vmLaAdRiY3n/d2rpqqLV0JMWAGJI7gPu5f5pXcGKl43tiZcos3
0emhxfiSyuxQ6lClGJxLN3A4P5HkStU0yDgnw5gobolbUiTJpXEReuzU/Nz6RMvDlV2A4btevFBT
7GH7O5s2dSiwCRnf5vc+VPLCaz5SZBqowg/Comp8I7H9Ms1DkyhWc9LgIIij2CsUVjOuctOs039B
wDjoLUtRFArJaeM8E1YIheK8xbdv+s5bEFhEYmwdC4o9vr4Ubc9u6KsxTAtwEtQ2++h8nQM38ZkL
sQ/TIbt4+w/Fcz9iLTmUGCfnPaNYdJnBPzgP1J0mF79g61geErKqcqHj60+ouWKYahUqcTRob2Gc
il/zcwKzDMHEQ+yDJ0IBJG7IrqMv3knURFBed12DHDjpkrcHEMGE4H5GzwSrwud65Q2z7yrcMT6u
KzgBd4KlMaTJOTnCOy26xqRbMcKN79ewjSsKyLmUV2J3y/lkdOZWKfkXFRJST1DA1r6aYO5jcZsI
RxKHZrekBAj0fLFliYQz7+lvLalrsNwjgKP8y/3VCOTiKbGzMHJ1ZIYj3PJ7Uf/eyDeW5QQ0xnMT
HjCegwy9ucdEn9IEJF/h17u9Q8VLze168jX7pIFGFazY++kuZvqx0WrUX1A5D2F5ejQwOq4vgGT6
4ydkf0RIb0cjMFn3/ibxuyaKF1tLaD903aXhRZDn5+s+Em6oDlHij09Jg4Y21Y1lqTW8wmiQcGuO
q5MF20GxVjW4EP09QzujdZd1mWfYZXY/CtYkJN//7ZvqLfsbRiF7e1Rt34l7/8K6RGCg4ap5FQT/
mZ25ZWpqQjPOLuMPRkLd9mysgjIOd0D0mubyb1OO8imODjzblctR1lGbE2Ne3z1RETJPCIyYjsTA
ay9vR3qquE63Rild3g3lfCGnC3xgpbZm9C/xunEdS9Al2nV0A3tzSwkDP0tFwlPTwZRvLa4+PJWG
5tQYFA0H1dIfJbMqjfy2b65VFswWMLjp1bXGJZRlcmogmhi6jJYhfCq0TadiBhQMKHycbxWVjeUk
0/hxgss9/xYsb9ihOkK6dfYpqOwBFubZr6X7RP/MzPsc5yr73Bm+g+5d+Vv4YYPkPDOdfQOFX2Yk
WGqFLkaIix9GQRXkPT5WFjQ9uMM9C8AFP7i22tbhEUuMKTseTdfrtd3G+lRscedbbIOoXjGTSHcQ
uH/wzPAExONDmi9XS/4pRz0RdwylBPsLVOaTxowXqJLdDfYUMaviuCgIyvIZO8/u+6cG5Vzz6VKy
RnpejN7JfG76m17DKToqUQH7GPDyBsyvYH5Z/tj/NRDTEF7J3pOz4/fS73x9ymoK07nR9qzMjIUa
y+J/yxNcyoi5TLuYhsfaJJTNKLRaLw05Q5JAtaka15y7M/pVYCZtANZRMySd//Woi/NmcnKtzPGV
tJ9LAfADKnDqJ+RxGcuY1Orq+e2RuU2bv7FMZIwkdMdu3iRn/58hhYyLCnKeO92giSQM/OBZEJ7w
AdrHbxMqTsTgQ8HB0JHym0Wet1FxnLbIsy0FF5eptU7XHuG+xqdATE3vGSC8JTVOzDJZK9kRf5I7
vK5e4EvrOrDC4frhlH8Qy0dWJC70gUUn+J20wz1j+72NX8GuA/iM6p3SUMPiCmvry9ALeZT4RvL4
Q33+kL4JCU75t64cyREsnW4riLb/jcm8aD6qWad47TUA87u0SBscRbPmnroaqzfvS4udH9v+xmby
XdLeI60ohgOhCGU/uRUsI1L8nzOgRqQNccOMoh9eEKznUfvn5haNnfqNE7T8Y1w2xXT+/OI9S5e2
tecHKZsdKDDPjYd2Mm9JHE/LeBsKSWDBBWY/BB3cxk/4C7OlgzCbm6E46Oi4ypenPqL9FYYWh5ES
gTlGmcwOdyUcWrWUXwDu9BHS/XoVPAE16F9XYJO68kJNpIiAIEw/ySrVH5vBQelkrOnvQnaLgZaQ
HN/icXvKCzAx7Ici9iopj4oK0s4W1gSjb8P+7riLaiiI3YIV3n8YjCwOODfEOQPelxDC6hQQlwJm
mQIMUBnCFPWp+IC19J35Kkt3pnHD5xg3AGALMPSE9a77W0SOUxnUk7U6daE2fp2hj/+o+ulYNRQI
DLv2NcO5LrkWKfmrAW6PjwN9110ey+2LZIX28ijIDkDp8xFeAUOlkdf22fIRcs2CrWwa59zqIBdd
yJt1eCds1Ix7W0EmT4Ca9T1YjA468I+fjDkB9QXYrs9mDhP1UCsZiDDK0N2Hl8BB+MsBN7n9lvug
739rfKNeICAn7jdIJ5uPkL9rdhPYnxsvQ1tBnl5oz43W+ILpL5e1qP+F4ymNh9ZRe0ZxbecB3s46
fCbDM49sgORwSPu+PNxmEl7UiTg/b6sqPV0eAsLVmzvDyPnWQasp9KEObtp0McdArEZhHrgd1++v
X0VYWBbJVbWmCQgUX9SXCJBdRQ3kVBBZB++wrdMSp9JEzN9wK13r0OkrjAYWj8kOKftmP2ZHe+e8
GhcRLcAx5a59fub2utvgZJWsqFy/XC1fNRedOIGUxufxUtG7wl41ZM8SVACTTXhQ4ST5uSnquS4f
oSd9qT9BO7ie0Mh7eXz3i7DtZH+DANTKSCVZOz237r39x2vPMbGQYqSSTROhx+gQyFsYeonoS/6w
p5WVE+cBg9hxEcfs8LSh3m84KutAEi0v+zlrKRDgstlEZkE55+UUuXdXvq1DA9Amy9vNlI0X5AmS
S7pCHVrUAZyQlIdMoHG5/VPsT4Ht0Mf2RK1TNUKBam45AqPKqntbqMSo4a9LnU1PSoCZcXC5E1qf
Ba2gspVCaVT65X0JpNnN2IGxEU24k6xo4VMRGh6tFIR2UiWKaTaoTxmFKxBFqBfAx0mg7viWi2of
NpdJQcNZUlQEUIyATy8byEEJpVUsnPxZprJxG3cGxHVsRpaHh6zhWvJ/FJFlAFd6pmtW8tY7kcJS
1sIn7rxyJBJBW7LxB4WtH/n0eTNz1tbtnTaGxPVSi7M0Nar/qoToSIC3cEU6vjkjm0vl3FvkpFTC
+taGSPQ/rxuUxPMFYUSHZd1RSgXrOd2HfzbTnWUlrddZrhRTpJzKhmB97TSnZaLV5nQb+prXFilF
JY5AE2KG5lQc1OO4xyu69qoUVFVHYINeDeUClTU9rhcNtqjvvv6AFKVWsg0BXHduHD909cQHPsGs
TQmz+Ph5Q03Pbk7wAIsOXlvc723lx3TaqtBOcTo9s6GF5ABeAh4DNBs2zD/e3CeXRJyChwL8vC6j
V6RhrEz6Hd0IwKJh9aBxMraeWFWERaYM6PiRWBfxefFkFnG8KgyD+kRBDMXsJkCvMqSTIO1tJ4RE
ZTI5VKrQF95TDQaFeIV4Lxi/HXgiFcO/zI6OQkCyQIkhYbAkRQSbXDWEDxBsWgZop5nOC1/QG1Al
XThe+i2U+siKJrY3MtQP/hhXhLBM30ZQpITvv/YH35r0uRZTFp7O/pCK2kio2ajsXCCXsrgDSVkj
hwRjj01hFqSUgBVHcusXHXc0BuZ5oRursYHiG7pzwaoXVijZs8EG0kfYl7qNUAeGml8h9GUt6YB9
fP5F0fS5denx5LGTgG4xWUoKu4brZORbmb6nkdMi6STFdUpdQJEDnvwKp9lkt2M492CTLgOYklI1
Q2epJKsgbyz0xRJN52S9Lxb+paoqXn8hqbqWa28RJ3uKK4Df76At7imvZ5WPi5YmdTLwJ64CS75Y
zOrrjMQBd1t77l//en6RxEdpbZVsO1ztpw5n61A2vN5QU6MPF1wPN5XDVb//MnBzKPHr/C5afLKe
oNHOkCw2263URsnewIBqcVkZRfFBj9/6FjL/xPNHnjSx1x9la/2H+YX15cX3CvlS/4r7L7l9LqKl
elODORqTU24O7znVhzsZgur9Hu3NfjUSF2sHuxEUjebppeDhseeaVvs4bAI8xlnktWsZHYmRjSxI
qx4IYA3u09RnFSDgH5UF7WiaZgyaiElBgRgK7i1aNUSAdWPNcMy9HeTvrEvqiuD6lkpfWE3flSd6
MD1r0lnAWsCeACjhuafFQT2Uh2vlwGFNHlMu90kjAy/L2a5lN+T1m4Lfg77GR95TusVuGT9UMqlF
PfWIVUxB9Ku+Zbchizd3wM8KL+146xz+xkQ9u0QHVAA/MLFi/M9u0R9KIwQl3yKkX5B95TiTBNuE
eIJ2BRQx6y5CpzXbvtjt/+qpRMK8ZuHU1PbX8iOjt2XsriVXPg0KZY+VGmtXHI3zW3skCdzq1+ul
tlHdDibwjy/oMfBSljo1l1TGabw6SjEfL8RuOOvxLtJqoN7SKFONzGhyR5gn16kFB+qMRAYcwhfH
/wP7reKVwb9V3S1V3K88xwkKYdi6jr+kfisMz1nVwgVauZpCo2934KDYtLdY+JKKW1g37XwWzvH4
y42Buo+l3OTTlPw6N4u0RhRIhDN/Z2aMa1McqGlmN0bQOSkMMpaqcb+mT+QWWBzIMGV7RFgvRoGT
d+RSlHFrVhGtQAgVhGXMgsstap+4n7J3USHl36JlocQSZqvaiXoDJbNLD3c015gjVfoERE4tVeWf
z9LNtfCgzvE2TuN2oUmfPYYrMzTdAjWWtH9JNjFZ9Xcu2z6NUb8dehVLziDQK31I1Y32olT/1HC6
WnQc2YlqFwOHH382k6SHoMAbdgYqJFugXELAF2Uy1J8+V8YPbzesDUaS4/YYabwJkoJd8MOiOfNh
nDtnNn3SiccVCri385Vdbatfm1eSsqqelIDqVkoaPqDLu3um0w+dL2XtX87J+bhMuAj7TT+cahgF
jQQX8j78MgPzjFtkMjZE8CmyS455Mw52qHW/kKmpBMtVw+Tme8MkPufrvUB3PH2t2dOfVSA4xWaZ
1JLz77rDi1EKtcaVJ4jNMp55Wn3ch7aSmhw38+MPm1M/k4VubOSROc+ZIlvDELt0JH0Zm3rBqVQ1
d8NLvvwvKQ8Lhw+xfm7vF5sRZ4yUrpUdNZTnJzd2LVvVCa6IivBT9cUYDRO04umIqV2DluRQ7vnQ
loau01ndfpJlFjnPWUo90F2AHskKHFiLaiF6Qj3ex69REvMxW8l26f1aJD2snEvTKksYuQs62yTA
J2i71vibW9wW6KQE/npYXHMwfNNjSMv+XRVWTdMxO9B4fbp4ceAUPKWf1/Awez6E4xReX6BHlTzQ
gp+T6qW3bIpi0KApNpp2O+VkHJcUiO6CrJ+309YPeQF4dshOuY+x51wOdfjsfl1sdCvGHVYZyXv3
s0I39jvgxwOsW2h4GQXvFwh1GdB9OwtjhkzNMYmI+VGBotfm1taQSFSdhFEOamY+eGYRhNoItWd/
HvSO63Q68mUYlQbBnAgOGIyC8lYs3RH6PUjAU38iuKXuq901EwcI6h1IEPvgtrWNGSYhnmxZIm0+
m5v9KwYw7AfLLqswVMeoFfvjtS4y5XlUl0M2ibIEWUTrTDdUcUrQ+pQw3LeTmIF67xFGMha4OwxR
yT3N3c7bGkvZf8fD/fMtHsyvJJngwyNldZ+3xORVakMA2abPGIfynGYOZV8U7w6AvijiVes3T4KP
tC6eeQNgvyZd+mr8Bg8SO7LB7oJHSmsRShOv8SSQIWPkuwI0N8mvd8bl7FX473nUepesMp66Tdc+
KmrpC7g4/B1MTMpbRzuJ/gbx+mFlIU55O0QH0p+BKjxl1okrLp7SN+0ggB5PhM9sC8SefaXu45Gp
HIe5TJhbOIk+COR/Nl40lJo+TNfxlyu41B22gvpuOYJKrAfx9iKdVMNtEIC5Jo3iq4DY4ExFShf4
hyzi9VpAZs0TUO33FzjwYvergKbD+nhwR3mjJPwBxTGApPSoU4sVLHVdOG28ZFOJk7W7DaCvFKsu
tGF0Ng/s3L6xABzkg7IrgollWBi4nOWcQD1NTFlIK7CyNvpAUnYRTEtf4Wp8iQMPUot//+pHuaoR
wRjTLZaR9rrqNeuWoxrnQk8gUohVvph7i09imICK32WuZ4Wh830ATulV8XACI2MGfgzQPPR1nZ/o
bj6xZMz8wOTjQa+jEOmfCBwmTuvHA1HzuCkBYzrzJiTs/VQzQeACk7MpXhqbk9VR3qvtyUrTz7OJ
00PyyJng7WuMd8t5Q2dh7WfarJzt3D4R1VdD4bPG0moxLohJIFT5mEG4xG4j0mhli3vETr1UgONJ
bJDJKcgIMURQQ/jCItPbbEqZUjIbH8lu6i8OT8m+bVS+O5mXcFCPxLue/+X3JZ1DcF9jtcgLJeI2
SDo/xp8QjmcjZiD8IlgVyrSuulGkcZblGNeQ/pfIm0FlHn8y9Mnr6mkHfhsIawHvsbw9O/9Nkmd+
dYb8zYHi2QnkrDK9wC5jMbFlXslDdmH6EyhFuC8CS3v3iY0xvb4tX3cKnIyFTaj86UD3sB5T+AaV
pNcK4v2WO1OPCdOUFSigFyWnqQT/FxOrtfIF/EZdpPcfKqgTDdPw3VqbaDYFamFwAna1qVyRznXy
aEIUp2qUvFxGpFhnjW0IYtAZyP2tDgSiEfk3dBeauZhn+Us8KjaHacZYBxk5B9aaY326hejwL+fD
XbsiCICd0C7YjLV4g0mRUTgbMo8q8n61tF+JJFJ1EITDa61s6ssdxxjwixb1crnQtfFcc1spQRS5
pdLTWmmU+OaVf9ddKhIaKvBeVDNrS9Fax0J2n1WSVzPyixyU6BJ6UQtkLy7V5cU8njagq8uVKMkF
kn9/RV8zXVHGcB8yRzCfl1vE1mvB55yeJFWi14btzX9JivGD+ZPmxu3BTsw4m9U3gxVvtn3piBI7
iqIU10myUDqcKCzlxM8IKUl5NDkfWPmz79nGp483ihoUw7eC5AOfsfKvGJIR5BBx4HLSagTTFgh4
FaAvAXAG7DgUAvPtSQ9rTvZx2F6OyQNk5NPmJGuhwJDCiGJEVcVSferHbgpC82RV2YPQlH0K0atJ
4JapJ02JDluVZbhObIWupR1XvIElh5bDQkaHT9cSqFHGnarn0HPurKiJMzoXHMIq5WGjy2NI+vQW
zmAroPpp9oJ3kXbHsIHzCppPZxQ7Q9CuEQFlhO6p0f138E1efvclcP46WznQYbD411bDCbS/0Ois
waRhAkVAYrTISN1WYCqt2p6gbcv08w9QEBlLUdHyKs3rProO5CXs1uMLrMkG7DfwOOGpdJ/lxCmP
ayF5VST7/IMG1sRPRa2Ee7lC3YUQko3mkuJoWrx2V1PMI8KDNOSlH+8sAQWlWflN7vdTmcdsbyuT
dXhsM6DUlFbSweSpcNn7YlU5zYQ3f8pPeg0ypyKGUUQ1sZf1uMciOT7+FyeLYFYc6Q+rEE35lD9q
UEHp/VNixgcfk4MvDjPCpD2iyM+GDbQbWnvbUCuOQqTwP/f5mXEFW0xkZzbVuVvw3nmN2U+BjKa3
YpgvUG908T62+bLm1YQLEY31bcCR09bnq811qzLQk9e9AwFs/9C6d14F4pQK8EGJ89FlqlFSelOD
URENbX9SLU0sr84OdkVALPTuI9zq1GnG9XJWKRc7LgcuCrvLlX0lmvQYCpAgaH9RM1xcZpjP6IAX
N9Ck+K67iBCzGAccEaMGLq8IaCZUTNXagVlXDUPyybKE5PxsmSuUCkdZqKbDfc8TRdKvCwZzbu6d
lxkiL3bRLxwiBNacIrkuKMxzdDAFDB62bP9rM2/fmxEn6vuL3s0GSezoV5aOTSrrPzi3e/owTT9j
MvQZV95xmM4JQ6QFgxYbZt1SvE8nUPf7WTzK44hPqoIDUXG+TW6r/kWHVHxt9Tjk1Q3XQaNBMMJP
pkjcOhiQG+r1WO/thzAY/xqu3yyQFnExXe4Ub4z68evHBXVWI3boHj50gQhkGJq11QLB8M9ORuH3
xygpzpAxtwNxaPVu+qWBa9UMFelyjg9XA7pu4Q2WkVaUBr6rXsXP46Nj285N4zh0LkrpJQjP3cz3
dpiiJcN1wP7+OO9Yp9vPIDSvgGUNjx6z++ybrIG2C+mgGa3r8oUFSzIOaWPaKpNgtuFoYn+XXCVL
rmtau8znxcnLc1kPFAJxYF7mmwCr1kE7jHCbWSrOitcQOpDJh6kRqNf5/UyxQp9iGiRQ82pmLPmK
6FC8MkHiKjDY9If8LmAESreC/QF88qgZQBA+qUgkRSzXgmck6Q3nb+Z+Mj3w6doaAWb5eNvGhfIr
oC++fgZPCkMuVWKK7GV0/rubKDIWIR+zFwqdZJrbNrjBbgwxiKJtIGm67808SjEtvBtbF0vnB6mp
kwjR5+fqPWZANNclHsxAAR8pgW1XeSevlm85lkQDF6DO+MPASM5KjnC4P4PtKXPu+8GDTRHFSY+Q
OHPp/GC9S6vNitEq7TnY2rSAxhZcn4/BUb02BeEvOoTRoTR9mtAetAWR/aPBP50j0RdKBi9daIkI
nI8Yy1Gk8s1Oz6UN08IQj/Hlnj8BSiF7gEgUKiU5xbhVV0SLpRASUW+Ne1Ef5mEDoammpeKHLu8i
PhzsEsfKAPAEw0j8L58N7usgC2IMRfw2GMHqC/b1qyR671cuZr4rIJeXNUxD0U9CrWNo5y8hMI7e
gyAvSULS+Pg3ywBOtPC5TKjzJd9BfH/8/LhEdypRx79YsJ2Tc/dRkqdqbcuSesp0a70UrX7toX5w
YRQr6+1Sain2xTH2BJPXQgI2Q2dyznug883nWmXGzf7V+kIEn+eo0Se/Pn/P7amW6GHs4NtBn3fE
OwAqEWeRS4pdd5ADoorqA+JdqQGAWlMnR9fEGLcrwmPsZ516utGrdPxfkZnc63fdVZ0ce4Mm5+h4
SoUxY+ETLd5pJJdmWvLvX/YAhHmeLlocUNyke74G8fc1O2NAXKP7dHYvMi+FjKi4rqfE5xeaVchT
N0PnN2rSzmgREwj6Y4zUGQw/7wOsXqYe1dCO0d0usgiieqJqDsoo1dbG5lCuVx3ryILpYS7d38JN
Sd621DlGNARCsuhMbH3OHTmKDlABb5MVYhgEihp784hI/frk8ilzfp0J9sYzm7x3XHwlV3W9kgkz
A7DUosS8u2RWGg1/M+C3WnzUGDP61jASiBD2Rul2qYVStqKRY8oPbG4stA58BN/9FWDCFn7cyK5C
22+Q4+ckl3jfcIGtzn5CiJkTdMLltrptEVyPWL1OTCcP/gLyylWovkQSXxYz75ggQzCAblw/84EP
nZk/z+k//7SOWm5hJ0AIRdiMmKGT1UrV3sPSvKLBzlPM3k+9DiEfceyTkDwELGo/45OS1eOwe2sn
mgiJPAQFCCWemBU2BeeysRK67PU5CZHQFiuBBpCBaOEo2ywvpE9UxEZol7uRVZu6hsJ+Xi1Z3lan
pHhjbHsNvFa2BPSOc2+Cne2+DxcgGnls3sev9HK+owHliN0t3ZjchK+1R54cSI1F6ZK8QUfYRJEF
4sDv9bXt6qBoaJqgRd1XRg1JJVeKqv/zRk8476/EEY7c3WFzJg/ap5QGRtec49ZmK0XlQGJ9BBpu
3P95zb5dRYeTi5VH09qJ2yZDc5gy6QwDZMCqG9UWKiplDVzWbLdv3oIi8aG5QI/e1A1GELNwpt4E
nyB/x7BCdFsZ/u5P3dZzkTcojnBAUbdEyg1EO4T46H6rj9VhJRL6DMMgUou727I2jxpz3ZgS5LMu
hZPux+8TMiwKUpfMXdHN7WRq+XHXpR8BvLI3nQRWr1umhQJyPWRlU0ylWawMbUzhbkY59boxaNaF
jut2O5cnPeN143OWry+2hrHZG7kxmoAUk9FGv4PKTB98MpLjoFEXmGm78+xL+lKzHc31xPyI1Ruf
loXis8B4+vVbiCDnn51Js+FvI4uP/700iv0adj+MWF+KpWpl+kwC2vTj13Tu2e9Bn/rDAPL87pqD
K/mx817IltxZfc2KFVYeHsNFJm/SSrORA15CWNXLTLtlfjow9v6yMAeV3h5NnbE9796TXEzjGnlu
Mh6tg5xDncG4O0ArgXzLoBe84JZOTJdVOItBvyR+tsgryFF8IiUC2BFd4VvR0G66k1PzZ+lAlHkV
lza2OoOMTG7T9zoPOOFCe23VnUxpf0DtyBgyCOnobRYaCjwGQ2PQ2YoVfVG1thkcaa7R8Ur8D063
7DQSkmKDKb8TJXfVelOFxD5vn0r8Acrqtwjgn16F/LH0ryS09YNsmQe9fGNt3bQdQi6t5jQgyJf9
5AfruvxCSkQR74Fch7ueKTqMaNrcCa6MZsQ+3eZY/+zjF8bYtCzKN542LGwyZF+0b+M8Qy9AuHvZ
9K1bAPx9/cjNNXoRYOvFkVOHkMU/OkbDXhPoCw3bqS1iVY6obDN/8eBO9AdUpXO3mPZNhua2v39x
X4yDZqmRLiIMBjnnDIJF2+buuRyF8J5QlwLl1Z+iqHIEAiVK0q5+hKqUtBXIWi1ckrMFsRuA8w38
1HM7X4LVpcjmqcSzk2huSKOlpJ2me9jcwjIHAGDaOTkw1pQd9nj+YoVLKOux5ZjqgoIxZj0i49BC
dZihq8vcPfFcAD4BAd9u7bM+uBRF1S6w8eXFo2v5n6FQUHglj9SRAZKScDh8M+Td1faODubq5TRv
mzNfLJ+Jm0x0SSXuWKjUNh5OnmQwyB268FSEYwSy+7L8k/CC1bKLJZC6hGfOPUFqnpo3actsdRXv
bZw4xH5Wa0c0qI/b+I1stRe66NmXi95/XHgJEjsw32c2I0HPxAaJjz42rMNhVtqi5ekbpe2x1IU0
5/xQ+ybYMEfTqFfakE5Z0OzSuV6ScjMiv/y1/BnMVX6D58++R7fOgFrMx5ljYhgar9+JGVYjMveC
pCbZ2MBXni4lCZRoPWv/Em9QfEDSZ6UZx+hNtrbvkgQSNwTx9hMQU5dkh36nUiGIOcFSAO03q+kB
O4O3JZmIEbMp4GKpMTsJFzzBekgIh4m3eV2maIONBlBUBEVYFYSNubY17xE61c6IED0RqYs90UCp
UkqKdNiL98WchttkipuP1iwv4KS+qTIVTjrGXnF8LPGIEddUOxHUPqi0SIVTmSHzQdC7yNLx5CHd
YwNb4z9r/DH0NpPA3mABA9dCbgSIXBWjp06P2ajkED4NcIfHuU5npNcEX1ea2T3Yce/a+REI3DF3
RMOrKabdUy7xIzbwdFLvFOZqyXq0h/GcsafxFDyJxOfpXigjMMeJsaoKmg0Pfn6fiMkqR5D9f605
lWRsg+w0MYh0oJ79OZMqXcY5BcwyHxPFDHp7WPpwjdM6N6o9qEFsAO8vwnU7amWU86Vz5GqA5jwE
+1jdnAaY/tAVb3naKwON2fLd4I+cE9gWZgnSHqw2xH2eYcaOHE/vUOZfyw1jJeb9gPgiB5ahFqp4
TIURY2avP2i41H+Tfm1m9jWHWYbUfhzoq9fYbek4nsIclwRwpy//lI/axDxTnCy70DXQiTxKLQ63
QodIH2XoQhbg+iQthw3AG7gjIiiYj4Anj8AErWzwlyhTwJpX0EsW05I8M9mVz7/vSPJ9x4DWy/KD
LUBATGys8xLKz+lZCr1ns9O+NGWvK5V24bJpJZbkczViIVG7KDmMgtSYCglEgk712rh2AJq/Iy5I
H0WdjWLBb5Hwr8XyV4y131vjmS5MPpiTyv7Qw2fvfxtbORm/cST905BODAAyl7DDtqkIcc/bCLeu
I4Cx9AzzBlnLuW2PEegVA5LHdgg1ViGPSHrvgx6KwAmno3BzdI7M33NAq3BKTeET+HWUMyI1xV1u
VBcIjYWvJvcWO3v9T5RBJWGLLRpccIaRVX4w5CCsCMyz/I7pjEOyar15DqboJ74zuLb446D1o2zF
UgbDK0yF5qZKkRrVNZfCsvIPirE9RQ8JY15/lwK7Jbz7joG7Y7T6dbENfeR53enx5jb1mDXV0mZv
CTiydn0ds02v2Npgr47uLZS5bbADHYwDt1YRrvx4gvwuyn7/FI7JRtF0yNr0XFixsY6pDiz59UvS
gnNj5R6Uv/Vh4wTv7Hki65u8oU5F60486x/dPUclppcCv17x9qF/0ZeA0nSDA5G/giFkQE6GVdaw
fjnjCv0qrJ623rtaeMVYr8pgbZtDrWKhluNUnA5F4WZ41KbUvDdZ2zSQ97FWjY6FFaugMzraU/UX
C9g00lflPN6DE8hbkxRquPvbxlzqAMM6XPjZUXp2HkQ4IPDdGyb1Sec2qEzbbsB1ultWo1iBwKxd
cOMWf/TUt8OTws122rj6F4j+xS1oQE/rbp/Yb4duVWnVq1KpvKyXAqnPD3PsBJ5JKsY6LdAWaG4e
MtMxoHfmonD6VCrsFEc8c5GhaCYXI+Vy7vqgVCrbo3Fw45b9SAc7CG6Q0LUXMm4Ob0vPIEZDIrE8
ONnXYbG4s5yWIrEjY81zXcfKX7hSrnqAqA/FGP7NRzfb+ahF2qde17X7IFx43Y8rtZnY5Axo50KW
Iq1+o+3VlIz8d/+xS/BPlD8aunneHFRvzNdIIr0GWsUIRAffBV07hHitqhc+ns+b7k6JfUeUUCiO
LwGqA6N8n3F4z8JZcjnIANP5bPhQUcwuVtljSn1OxWwU7ccTaNIrJIdn7PYbziQBijiD7oOXYj6R
F1NphhDw854PwzWJxcfzh4Pl6DC3KWzWR5O7S7kub8EAtB2JzVsTwJk4FFO0P9DHY76JjKQNoleA
cKi/KMjUXgLzGA1exaBk5NlTzOVezH0jCrKLjyihpra8+4f0TTecF6wFlZtcS70vAm3EqnC3cqv2
VxfTuDzSNL7p2MJ8nqfFz0uojPNgW1YWOGLJb1L9Yh1SNZgHofLoTWw2VRH6P7eN6b4MKLwu3pCD
f/jSTOsjcegvscR5HVIaWvqvfPU25swlNmydBnQ6ixXg3Ytmq2D57CRJXBqyTh2u6XJ54gqpv9Fl
unigqkk8VamMB25q7WIk6KMAdWGpwcunQk73LzCdQq/qz33ejKmgf7noNCC6VbZN3hHP+JyskhK3
EkILQoZpX0B7lBjP6OhTmrctosbfCMD/oKevzninFxYMp1PtPEAafXw7lJbZZA90AqJ0Y+I/SGBA
9h1KHj+dT8TOzPjCQpngqiTqN7ZrOeS1C7+P624rIBLF4ZnFd/O/ynWquCjRzpH0gm0+mskFbEF/
Qaps7MSbL6tOd5c4Ph38n2zowPLsX97N+Zf6xk4r1ItKhwQGPC1p/QlTNBqPRw+ChJNyt/Tjt0hM
nLYUpdpIy6rnUoQfMzqnAYSOTAuK6M9YFEhBBsCZaRBHuGws3HgP0AKV6p86iSvOxsV71GcdS1gY
KUr030szxiT5N84W5W4Jdx3MxOKpDqikPVtL83CPB6LRYhPXvo61lOc012lmvawCfxko/vX//DPK
1qCpuhd70mF+kYABbVIfsoxW5Eh9SjvGKUnmZIdDD4u+ZKAa9JLP/seX0ra4WTqoWzX7wav9ZBC9
xDUB9bWq3ffuxD1yIGRE7xWqb5hGoBlMddGIoZouAqPNTvduQIs0upsQsLRV9/gqzWe7u8n4fPcZ
dgHutttnJI1p+aP5iACzV3y29VP7Y2XMaJx1MkX7FrrPDEioVg5BP8BFE5ZdLZCt6ShnMX83QJQR
byYPwKd0xvKf9Ed4MKnO/nmIAsgfedBoOQQcGXehD6yCT4RJYw/5w6y6lSuXGiWBZcBcauAHUjcQ
/5mgu6tvREsmPMiuxg4n2Hdhjn450OryiVwIGAf0arX/cFrNkfidlwraT2JgI+aUnaY+3ZVuSomO
BIFvL/NHJkg4H+z0DixV3J0V5dNxAQ/ZNXB69tG0+7DNmunTldYiTbZ2sAa7bGkgbwm/h512sfvJ
ffDjTv8sf6l9Q6mb4IwB5n8VxbbaSsRCHZHbNmtxTJ9lUxEyTc1RBCciFaiCzecPzVp7C+9FjpLM
jYZP4tW7Cbx/so75BRPflfJ78zIeIDKEwX3URQtwDfjubEMUBiDJJJanjiXMHjxAdI8HokjCMmp0
1AUb83QToPM5PcYRSQHyaJB9M54PbXeIBQ3YZ84ILuycWJ3UR8r34XhCU0qyrQYU9ATCZT9tf3tY
Dnr2K+eIus77lFR+6XwR36QTWvdUbLw0KWaG38PrANrPXd781PyeXeMrdcS2IBSkArbBHf2E+vQc
6kNlBMuMsy5HgoXlrSVCNcijSpx6a6SE4/o03lTq4xOnATYZvrOYtT9SLEvEH/+RaFzKJPJcT3G/
FS8xXqQg96gCvdTj521PCp5D0ovXPWVntUoRz/BrJfZFCHeL5dZJr2J39qx3EiDu9zjG2kgVJMga
Mw1ottCdCwJSv+SUxknGYvzRbTUvSw42AUINio35SvqlySSY6ezaalS7iyyXdn1QVEGsaoJcB0IC
wnA1Z5uC1TClBQ25fHkZ6GFbPQMMCCeCc+RK4Vi0RlRMnD6otWcV424TDCbRTy+CJcxqiGhzq/qd
a4f+k1XAl9pCg8gbVaMy+t2QZm2HPoeu1MBCBNVPSh87LbE+Ms7ecew2UQHximjpdSuMnvcUypLA
KoVPx0oMyd0nXwVqIsaosm/j7b0d3uImcDKrdgyVoYjvSEh0m5jTDhgPSZ4K5+u3ivmvKrZtoFnh
OGZrmvHM+s0YrFll7Nly1weKBnh91a65U9qqhHMOMkFD69YI2U52Lv74VrZASMb9gM4NvTvXQMY9
ULYZy4LAERBXbm8vpY6faR6szmLQDRmP++ie8gpkVxoanntHkMo6x/zfNjFjTkHQJ8cGnE1XQ6jc
23+rmB2uo8fZ5Q29bgqwq2PBFliXe4ey675p7wBQg9j0HppugXHLDyocmog2je8fcRT7gYTSKcx9
ia8L2shlk7iPbM+pfiVv5QWuckKt816LbhWXuRTj+9U8wSFIy2hF+3gqMz4nkac8BsDR2wgoBKIR
Em0e8EkhJySqCtvahzf7bNUjWBTsmBIBFvueEV0t3IdbYvgT+KflBL2Z+D/CMfZDa4tdrBoKfxvl
LL6gG+ElPL6OqFT1HZ51JNHdA8pXPvhhRqW/Y/PPAqMpC+Gv80EAeVcKQGDN7H77BbQZLlLraSyg
X6NON0jVHzWa4dlg9B7eRUbwR1kE+2OU5VZlfGbUUX1ozA82MWH8qSotC7oeFC6P3B0W11J38fs4
ztIKLiI2p643dIhL+YY45kspnmRimT6q43rsz42T3AHFaXaR3e4aIwLJHYqKgFN682v1zZJOLJKn
aOESrwfA96lK8Oyr0tGMG7XFY0azi0i0IdKmQT/SdgPYTSimoLl5dwzJtspBP5i3Kua1p8QB5www
yIJUUmItPsfmXWL5cIUrEfG0pbd7Ya0uVFZIO6ti3VWXDowSMSJKLkRui40tRXZAqCX/EdsmarFc
sato7UW33lz0fTDXv18Z7g9iMufWH+yVMOyfXGSoq/sWOG2E7VG6Gv+Nlio6L67sLBZ4BUDjWz4S
xgi3FTUEiO8+bIrFZL5hm+EcKr05Vj0A6PSj+maVKaO7PXtk1suePJHH5c0GCnOCuxsq0wswQen7
gp0gODMa85ZeZ657+3wkQEYGcWpFGzpJV2YZNmfbEjVVwuLttJjX+3sc4wSwZPmmtwaLw/ljUQRX
IKJ4fpYYINCIHNUstLWPMlNDRD3WOFQEMjIKgjECPL7sJ9qotyEI0V0KcqLxdlCkzlxbMmVm9WPa
fgjo2lc3CKdAmx1uDIPp6tpWySNpHOAW7+BPoPnJproLyyxjoGps7UHbj7xfjGcoel1HmHXr/k/v
Jkf050BThyffS7OOETqaW/OZWcqECzq8rzGPN/t0dN+e7gjbinETKoCRRYip5KvGFGMyEVscG4/N
n1ls3+/Xd6dmNO1kofmnt63cSVGGrnJKjTUb7fw6MjUFbDfnxtbfIxVSSEtwE/s5XFpqCPVaEV9y
0uYzaw3sSmu+1MqM1Q62DYvesznEMhwOzeC5qB4YKGn7/lo1udA4EbbOaL1hbKVFwQPnEflUQg6B
MDpSg9w0xIs2/njbiPiykPDXhi1cxDR6ctxWlq8foAL8aUN08fQW75apO93BcRkDJktibFTWiXNX
zN5bNLy99IJChC8vv28rmLO+KK0bvmiNISK9bJaRQA8VRwmVRuzZbcYNGOva6ZrAnIxfSuilCm4J
b9KmyxguN4HvhVcksoHAg2601ArwMxRhWwh9nA4jfN/6PDVH8iWFdGdqpspOcrzke7VNeCDt/D+j
NL/ThvG3XDK3sQk/22iEs06tdouIeVclcN6sildc/TWmQtQinGLFHQJFteyo1DHyjKtzw9Yhgqkh
xBeyXjk2xHC3ZvwXDa9XKKNjktXopx550uvCq5W2mChin3XyL8LMkHaMbBnWFZcxjSUZZ/sPRbnx
gMTvsmBSs0UWm0ECRotMUUN+7FNYZiSvxtdpjjIrkxlP3W5DrBRXWib26tDUf4Ce3g7ovyK0KGNC
Rsb6NayOGKptcGNYIXAfVolyXtmjbgrySrZccJ5aqXhr+HylkFZocbU209d95CJb/R5fwU4nlbxy
/TAo4fFJMumXBoUuNxKehFgg22Fr6Gra3ayjZVBBuAr3Ry0ELXfJ1yJfnMtao7SiKseTRCJ6TrWq
/NJ5+GQxnOUCWjE0p2SV7c63mM+bni/I5WbyhUXrXIaqgtlL9RTi5UByrmkPHKzhKMW5/IJmDT42
ZGOw00CItsi2p8Dre8IggJzpZpM0LTN+K1fuWoNn5SWmU2hLTOCPuT+BMrWDLXD16g6ROjAZ9Rxw
kTrkodfPYocHhXNsC1NQ45ZnyWrhdKcG5ILQe5Dwd7EaAakfWyIInw7jst1ofcrZzUv5TIQ7PN2n
FAG5Q9L+cIl4qd4zPdBtKPv1Fg/H8W02ckJAvHcjMk/TpL/z7oeLDBGM/73nJUOADtAcijzhtIIh
z30usrqSElWCfhFcFT/KPzn1mnCFMTxGaQ9DP9NVjWDyDDIWLADgIaN1llRvm8ET2AI2rZhR5udn
0buV44WhfouiGGLBGyPl16uBeNXey6Hjjt+1PwDcJcH6rAQ/AuWnmpzl41SgbS89IkKX21RY5T9W
4UittOolbshcDq3Llcnqq2UlK/12AcV437IhEOIqaSSELR+Ss5UM9yrzQinZxOXG8jONrYeAc38J
BZgXqyG9b10rndm6sHGQmL7+pgdwvXVh6K1rfoPk74nM95Hf5yudNSsizp41Pt65sTqJq9yyH7f3
P03keB3YCnJ8xWUrM7b+JjnyZFNSt6jrQEqYLDtxPLXsevE6ntrP3VIFJ/YUAiP53Oct70sOsOzw
XEtvBCGpGfL6fggs5x8inR3LNTMgn4fLVI9r+fzhzsfNhw2KVSc+Ny5EeEfpvWshs2ar+DvDdIu1
hU8LvMy8b3+EU9jHvpFB/pjH1mtWNRCgPEx+p6LJnTn9IzshaBXjfQA2I0P2clZzBZ34PrrVMqeh
OI0NmoK8vuebEFvmztlPhM9eSXFeKy7lwtOzyAlmclZcNhMBYZfRiuBc28UMK4EtyyRJqG0al9s4
q6PBxYPsAlz9WYKz/uXyTUZTyFAveuG/MN3CSlsjlgv/pNT9cZM6T/PVRKxXB5NHjLkEZgdZ4GOV
kSU5/6ruEHUn7Miv4enuSpE8njtpD54E2Pqx2r8W9PK/+gxfoQwiNlzQ/eqWOIstV6ZMFnu+eMjo
JcMEiY8QMjl/j9fOrc/SqmKKzPjAv29ihEAJT/QY+5xa7hmEvm3Y6Z4y5uDV9LQY6cEQhCActEOc
//dW4L+1iKPLsuUhYOXsudkPaDozwwAYOx+Fm+zGcq/gfn/xp59qAthq+zYskALoeu6thSMoYWRX
+WqcDNLRvyQMDtIbjocMeNrXVDhW4w3K1pNLVNCoEjYegZzoIpHkYC7qtIXoRHy8o/EGk3UNj0JW
eZKXUjJjMmLbuYxAy6plQy+xnxCKju0j+r+lKrgfJG1edNX/nJzXN08aNUNuG4qQ7uJ5l5lJPiVi
BPnW1KjaMxUJRavnCOPehvD2rWhCxMQUGVye42MsigJX6cdQPtv4QlsbrtiLtIBS48PY1HNfPE0r
SCxW3v5CqVcIdV7x16f7VFcEToduS0Ua5jtA38SRP6TGzTd07olFhDPoEdW7jwcqOUAlmEKLwU8Z
SjVhOQK3aPgzspoGVfr4tkqIBvLGa+wfAD+9lj9GHWWdvtnHQY5Q2DEoRUpidKgIqvoICUTZ6DJ6
jvtxmD5vcakcjsuJti6eBWqcz/yG+x3N+pvi9jOtR39YeZooFODv8/vvwEkI/7KIiHDqls7GRgRp
51VDVZpOBbBGap8TynI1koQPbbADI8kcO3RR1Tooo+y5sQDJMEy3Ea8sEH4SB/hVi4H7QlFlSZef
Ldl0acZzahmdpPSascIM2qMm76Axcg2MeM4uVFABHMdexWx2piGsBo3r9xv6sLwChDxFGVBHC0NL
hjc1aqZwnkbaFTBfawTIlSjDgN1DdvLyFnxUIeg403upLGUkdBxdjwLcyNZGw1BiWu5s47ZBihg7
zF27vIdP9/mOGuw1cRtYBnKnNnorYQdbQl2/XL+54Ag39LR52mMMWEEWTpi0akQ+pRWo+kxkGpXv
Ha8vBubQ2YAVQ+SQC0HE0/QvQ5AyS0KE6eVblJWjqPTyqv5TH1WPNPfoXvbwV5BrDXgF8P0HJfE8
ZW5/P43uQ4rAIEM6OzJvtC9wWRiSdZDUAreSQDCIQMEgsDJfXparTbcZnXve6oWpST2nixtn0k8K
mfcSVk2uRiEsS9o1k9F4E6IPF+7RZE2Mt0h1QpvEtSKKy7vEUsNpmJmQrSzDZot7nL20ZmCJDFtF
V639lA/MDEBGqkeYkUDhgh19IgV64yc4Wnba3qALx1nrt/GI2Doo/oWKvxxuLtZaAkUSoSkAillA
Dz0oQi0DSauZAChjhmB3TTUFcltvjRfTk9RxPX8VpIDgBIyC2EGmqQH2bsUmpGjSg2CGmpK9IjAa
lhhfQUR0aQam9XO+EqWJoL/hkN9W9D21Z5v/Nxhowwp//CRo/rLyBSRUDC0D8vTdnkg/J977WOXA
9ncPhQ41yXqCosoCqjpCTROtIN7I1gxVUxCfBau7i3sixdjpDte1js02cBu49Fhx54LZUlYNWRQ3
r+auaSZfsmhS0KEjaPDXgx/0KSNX57f2ZlazZ7BE63gY4DTrA7p+oUYMU1DU44BYRHO4BrnQ61zz
lcJhNb6V7qoO2NSs2a6VQf10qa9H2mkhu/f40qTNxwtwqarDK3g8y8sgE70KSaQphI0wH+7gBV4V
yG53mA+K7Outm7h/qUcB8skVgWWfj91XyWorLx1DN0thYJNpEVjcarucjFd8vtiUt6zE6ZYqTuwA
kKA2xqiPRpDF7BPo8hXascHfW0UD68ddWB5sPHtF4Mda6L5XgJsF31fcquZD95R7Y+AWymcTd6vF
Cj1eJc3W9Rcx1pi4La9Bd/1NAmuPOKl0brHwgqrLZVEkt2ZyxJaSkml9jeXRrSEKp9VjHzkeHA/c
Kw41xFi7w6Jmbo0GQRPq4KDwF6y/PJIWZ/kMuxyFHSoEE7xJClx/LQxfY+hZ1N9PrdDT51TErvVd
5P7bV2dHWx+ekogeMQbE6d5if7i4lxN71K7RJNTL7IZNimfdGaK9fNdFS4/SzEKXbrZ7Qp+lOV3n
KJAdo9FarVKQv23vlWpNckb11lugLVgzK7BvkPIpVSEqHpCd2XjzFD5Xbyf++Itup5+ni/ZNINqC
2ivueHKJryEWbIlJEsZly6JfXJoQhiVk1QvfglNvHI213oIOQ+PHZVIhSoplL1DSTziKytdYI8eN
lpsUrV0sBXw124PJXOrMwzgUKoHv5FABL5f96XSKItyjEwwMsEZJKNpdfT7n1HHi5Q6nIrse040c
mH6vPXgyDxy0sOHCQiYpzyp4BiV/nFoOHhW1fNoZIrmRc9gtuxgYOYl2LEffq1SJ5HgmdaCyMTVY
X0Hs4e3VQShFMcOefLMF1ApOxIhlHPpXabqIXvQLkISBNpFVMUN7h5OzWSpuA+y1SRuLPguJnAx3
YcEI5A7RezJKbXSMqFIYLgTk1ZCzLeNztW/D54AOioMmn5vwru8UFemu+1G/HhTHOby5Z2o5wN8h
RGIssWjLT7egek9Ezal20IdaCSZdlG+7MFvAD/INA6xBUGi1YY47IAs51IgZjAsmcIiWsKvg84zy
YvEs0yD58tRI7nv0vzwA0M353wJMFyB5amu+QjOmj3PZateUT4qVZaG1LvG3c/sH+78mazwphv/E
xEc8IKSJ3r2nANJzonKfwaVdQQOMzF35DLQ6qE7pDtdpZkdAKBqFle/1leApD5sb5ATzo9vT5WSV
5u7dTbGHGJQjDz9f5ZAOF5BysIAzk2n67nVVzBdTOYqfhpn0IJXutyhdi2bsulcs3XQ28YQA4KVs
ZScE59p4CBUpNKac/4JaZ2L5i2x96lXpsRfxL7B3cNbVfg+AiHZTGRmaoVlLV8o6cXRlFPKUXadV
OR55BfCYWQDLMdnkm02d7+sdjJHG39Jl46DFLi71nvlNHeCWsdhtuHwO79018IpscL/46VuUqT22
gXfj76ZfxyriK3gaD8ZVvoOEmZvgUUBBu3hdFNFiF+Z09cNQ93Ab/qj/LMyJKPcH6e1XDnOdAzMc
7c0xjBI9QpsUqqgV6Eb+Yh8/zNOEX7eJywzEcG+80gL6GIM13OGclHtSflTnMnajYdNDFGLEHDKz
scnYrza3YATUYSDVwKOQT96rxFCXYIG54FZBizWuPJhsAXFikGKyw/6nagQDKQiC/5cATwcICciU
mR2xHitt78pjvV6j5h0R9xzpvYkTJKk1AXPPHmZbUnfVwjE9wooJZX8xVaP4Q05mt1xylCSNNvte
b5Pec6ooofzy6k/e+yz5Ma7F4CE5g5NvdEbz0F1C2llTySibFqtoOJ96WzRL3s/Xos1LNlbiM3OV
z8x0wrV1tgFvzC7HiDH8saBHcgX0pNTc5dbrl8asA0C2yFRqEBXgN1o5bzYPeuxFRIj4hk5VH1zS
l82KRwFucApoW2PgIIsZZZCupbbD1sgfWQRstIxfnhUJQdGjl1xC49IaztdytOGx/WUmloOke7iZ
kDorCwODe0NKf8kygv6qi1kmCvzlRnzxztrm+PvfOR/YVVJQ5kqWn+gw6yVbnlGsIIcMfOMp7sEH
5MrHaqUpzw+fK7dxNk0H0ZdGLmFT1RlXyDYN6jD9Xq1PUdfYrLSDuFctgmUe3xwU2pX26Eq+WdYT
5goWDsaR/w/UbhhL3pINvdn/mGdu6SgVn413+Wg6Navf1+JcvUdIBBiSPzBjoyKLjW+6Chma7zqJ
hGxIfNyGdtF1s3zstjjnv3eqvscOs6Ra/304pKqqtXNO6Nhu8llocnwlxDfto1ZaJbk3jF6D3n2d
PaiwtQunCRp+RhgpP5fau879/I0LfyCJmmv+ybnY0XvoXnygipRJkbpj438Y9SHi1/VAzTqNX0U/
o+vlSVKr+y9ZF4jzBgw6lVGwP4rojVVd76A5zKPuFKy66d4wl9R0X0mwnQPFLwsUun9RYTBst+Po
jy9vywHcnb6l1Ip0J86SGxfuoo6xKclIBoXV0fwmohNFAjVUDhWs899kRk1v4932qAp/Mq7XDOFv
ZRVBBrcazrYrFJibHzH3G+tW5Xa7viJFCQ1pkCvgn15YNgdQdkDxegJMLMHSxStBWfklMA/6yahM
FgxOQrnEpy6XNew8uV7xBDTY6bPMMbj/nKPWxfzQf2XeGK04Nu52n9HLP8sdR/tD3cnS9I+HISEQ
AVcwl7zZjgj5c6FSVDBaJttiMQHxZxu7R9eZi8BHA8DGSpfrjgl2fPm1FtQmyMCopeQF6sDt+xeF
6OJZuTc72uK9i/9en1mT1c5oJLpy59JdxuwBXGtRvamj8v3zUDkNQPGzFVoHlDXHXjTLRuauts/P
mcU+kkBrEs6o5E23glPDW2F7ZrBL8TnGllX9s/3j0EQaVs0xH3iB3V7c7mHCs7yemraLvYoVwxVL
4+Gn/B7/WHtLRDsUAja0tsR8K4KCbawDATET7JRiu/d543Fy400uQ7yE1Wlv9TPWJN7JBhKzpGe9
ZUnUQC62bYHvANdbIN8PZ2itxqG//AzyvkFtLEnfhVNvV73MIm3V/nq6QjTqxT5+cisYEeI+mWOu
4MrmYLqZwCI7rgsoFtWSlaQBaXgO6OtHq7skkRCfhUNiI/6Znl7r5/D75r8dcJ1jWMdCYATl1qmH
igX9ixb2KF7TlI3ZAwUL/wsTjfcNEe0q97skhXftLY8tp99YTzv3sz95ZL3/Ng7kvgcToq0efac/
HC+vqtB4VlYHcBDpCfF+WnEFT7PLsT6rsv8Uo29p1ZpGaCfMS02MIrDeHsjLLt/0uVG4mrxPPkat
l7VNOIP66DJMUQt935S6wPdzRjxW8VZMUlSgoOPzP1UeGbDnl5kjK0Ko+qCdemrw6eT1+kxfNBiO
ETcm1udAXwQxDtdVmSO06wMQtOVT/P3+eeiWyNzHfDInEGoM8PjI7xehioFggGsRsF/jnKMPdfyh
84CA0eAvHfHi7xxg2wML8sNnmtS11HCFaaIC1zDkBoPtDzTGMjyz43kq4xRYFSjtCNW+QlaFgart
NriBQkpP9q4lwHUJdvmewjq1fWgbDoGWBiN7aGKSzpDLGPmea/BxfSI9WmiTACMqbQuMqV9W2+6v
8segADooRPyrj8cJ4FCGYnBxk9GfkHznug59albI6F0XuQzfyYrvUSnYs05rXAfv1nJmXEja96GC
zyvbN/bXx4001CYLoyzdKEX8wC/spVm53w7RI+c9Ichl1D1Ih+KwRsZ968piyTQTSH18rv9pYJYq
6I7geU2FLa3gWCJyjhSFo61YltuXV4KUZpGX7TMn8d0TBrilFuCpknUbjdR51ZBJIezPDosFGPLp
FnQnW7nxAwH723rJxGqHHUjNhZvpyKDushVPg2GPoTddowlPLp5QnckqTOfY+e0vDgwGtH7EUB94
2ZvWl2YD4W7Rb7Ic9M959DFbfHDPT8jQnLZw3AcxZ3bfzEVf8WzsjZBS5dvgE7Bv57bod+JdWCen
z96RP4yol/T/n4PJ2fKwjA/HUXSh5MG4LHfInM80rXxZPxXeyo+2xZwZPKuaHGDrK+flsuxkl/9Y
AfC3ble4/lEOIHibbzi82ATXoLPyZegXFcIXigdJC/TeqTxK5ig8kp7xkctRrfcThxARUxptQ4UQ
B5Dp9q83cQYL8DV1YqwW8FHrLQo6YrvuQ7nQksKKlNlVW+a6HJUl2GblmVqM6d32TZ8s5vfniXTQ
XqXWgZATeqQBkZc0vKtd92x+s17tdCphdJLZAR9AnWAolUP2FcZ/o3HhnsqORIzvW905qFx6vR95
prmoziCUrgkskgEWHKQkvigf2TapLtVts4u4Ej+yo6zAJc4vOMeiXUYvQtNNKgZ5sjDFSXtGeZeX
VyBGjlkUBruDAdnhHqwR1nZqLpyoiYpadjlXlROq1nXAWRaqOF8Vg2tAExNIp6vsKdHoggfkJoCf
XTofX8dFYaCfs3KFQHGEIAO1rTJkHL6jCZL9hKnWZ3R3vvrj1E19Won3da+s33UnGsUyyYDdoUpe
GobexSw+mcXIFeFR4+kx1DwKYjqGrokxvP2/G5AOZRqJSMlZRndDzDbsuYRqoPp1Ws6lTDJDLuQf
+eYex2hWClp4bIc5a0vWYl4E7JQB5K+iTJm5ysoZzp8GuDA9InoduMT5zY4/wmO52r6kTzqkzN46
bqGRRJDq61Q/OZkFQzbfJqhyTwCT58b0PCCOewBRFUszjYAs8cFc2XNWc/z6hfYNKuBR7SqNrWB5
LmmgEnK8jSDcRApJuPIPFg0hDQ2Pf2225ie1ayAeS48tLnu820stzs2ngqb7iovsQuk+DShcBl/w
q4j6fsAXH2RQkq6hX2C1BZuqLXuyKF3dCRm/YDXosDecTCWljZ3v/ApEwewBA+qlK8Xs/t3CoWVM
24ctEfNPBmwUOcqiC1accJGHW6ltMwJY+7SnEYmv2xws21CR0s6J92mGXAVKkfIkoLRVto2YUpap
mWoTu+RK5Q7625xp8RtdIvNxmGYYJaVR6Q0ZUwGHczuFl4fm1SkFYxMjunlqs4/pCVmYT6dySkk/
3/PSmkpAlFjltxYHyzNfKXHLH3jjbqGOvEOjHBM0mikTACScdOOAXO0zWiM5A8N6DoHvHUA48bRP
fxpGYOm1ze6QIIo6xsYktChLqt/il8g3npYzaBplGfLuNrl1P8LS54o8IbB27ra8f7XVFIkbyVfa
Zlsc8xoe04lDYSiiKI1NTYhCa8tA0kcQHph7VRn4+UA4/NPHNmptf2l5aEHStHdNwFk8XoC5BDRD
Y+E9PEP64uWAfP5kfojS46qNMiHW3i7hJOf1oSX+Dpx4if/9K4/AqUrLddtTInIoE/tsYHkqjQPK
MtSPvVBJ9b3x43IBCipjWTJtF4LyITTi/UAjPzzulWMH5cRc8ilPfeVtacmPZ1xwXZJMAz4TWZaj
xkPFKpJU9we8sxWpUPXGfOQr75J3Fa1U8xz7Hrl6ngfl+3ltvnRu8BwAKD5Eg6pwW7N6A03fYEkf
c2XsK1z29Q0lzh1JDk40h91UR3WJZ4PIULhP1kz5DBQ1JnOuWuJtZVnzU0fBQPUo9Q5P722sWLRx
zrNrp+3bR/Y52j4KYFhcB1azqwLoiNc19rdBOgEG7owH1TDM8mEyldwPiTB5sityTYWx2K8i9x2O
BXhK6xaW0+GvDRbs/1viK88Q6qnL7WV19twDM2oOlZzqL2JEZHUfwO9krb34F0Gux4ZMLBk3cFws
VDGCq32YZk7eKEQg3422voLWLCi7MR6wR0GR2Ot4tizi3fTBdDFsaXSMwUceRQsv67LqFrBbbxFm
7aGqhLO53se8Jbu29EuEN+qmD8WLhn7UfdGvCmXe2FrsHcB//UOMElTCjPbsEoiKcjMdsJWAJ/8S
3FyOI11zdnfg0iGTMEZDEzA/zQJAqE1OdXoLnAlyWFoprNzJtNOEL6kUBx6GPdwNCG/++MqVGllx
8rafFk6MoGUWWPQ/MDnWyeF57J/WqaimL6//cQElhiI81ZFio0cOl5Dljz8KvA1OUjg5TULk0uaO
/PGhl0J5Nkh45UKU6BtodL9JNvJituvNEBZrURzmjbBhdzmG10pmlUtWlPOuEg7A1fKXWgK0jdjp
4ImzrBHS4F1i5SI2p0Rd9I+4FoV7C8ZK3gdf7a/Ee6Cc4DYkeuPM9nb9WP8DCmDgAPh4+SrK4nQR
tWoESpkomwV5+OnJv8evhOSeYe+X3TmviLGgrUW5/fhRCYowyhonzGCwgRBCmZLZk/MN5hEyGT/W
QM0HxE9iWBZAINxJmyX2dvddUOi2pspT1oe3b1VGx8ViINHx3M3YkXdpagkft1Rm0zUqISTVJtAZ
LYfF/vXkQOoYEIiXJ560gpqPvLuQ1k7vcZ1hwwS0GWrHO6KzqaF3xwAxOqVWvbrGQoB1jNBd8V2g
gT5SdNAdbPZSDWTsdShsvOzM5ZG/mXFRv6uwumhHHiNe6/NoCw29veky1sP/9gizTEeRjzLvw5MM
1oJfYg0QTod50hlbBxCklPBq6q/gaiv5Pp/E2ID8RM3QuLR441Vrtu7lDeFKwAOKsgmXDSG890fJ
LoSeVUjjg5zY2TzO0k5rZWe7RiIXttxl5RbqQYQ/VymERzPktIXB6oKqbdDr9eqCsBhPxwKFKg1V
XHH9Js7rJEk2P1XElUy8cTQRobBa8GhLgP0Yw+bExQu43N/i6xB7F3rAkeGsSW/N9YO1IZ5F9Y/Z
hXfACEjkkUp3KVLcXIqE0x/OFuMtC2e972tgrAfkGlKuFe5pqyOJXXq0EhrSXdl/rSZf/gbMTDwG
E1Jx/eAK1uJq8gxcvGSTkGGqReG7uBvRrLqWw9+7Ji9tvM+ifFWRxSn0A6K+aHGBXMZljBFBoxwG
NzUW6rorCn5kEwATssWaf8jR3WpSry7sV9DDqpKa7B7b6Q2UgOnwHrgmeN9RYKOkqa6S+H0kme++
5Zel53u17arUeMzO38IHZiSMey3tLDhEsKwW7HDE0GvPNrf4+50vA28atZtIsEw+YWXtWYv5m+s/
ibJ/l7VPjg47tnxI/3qWzIC4L7W82/bcUcIwkz/Bs8TfTSwV78I2uAaBUTSrhiLy00SRXIqzWUiD
OWPqW+KlOmLKdCoaLSaAaGT405VjQWcCn/6DMMTW1nB1P98G7CrCcbFihm49ZYyvjRtxRx9vupBQ
pyHtIXzA1XRFXYjZfDlGxx65AOrQkPpzlRkD/ecdLR6W8M/wDMttga5RPlfQkCsdogJcbqAXftmW
obEGrqsZTyfGq6nKYlJWykV2GiYgO/bZShhAmpu6nVn1KYX2D4RBkHAGHENO2p8wU/liOVR6+zSW
BS03g4kYPBivVv9nuYM+pRCQCQtcrnsCVOkMRc5TIymtFXs6+BURzW6NnaRMNT/R1a0/WKZDV7fF
DY3FTBUuo7ALvia5oDIt8Wpe3n7amfewBKu4HtqJbFVaEZHmIMQB7Pys05XE2PLnODZGqN1YbhII
5MA4QXicQ23FHfUyJVuuouRBonDPE/Oup+us1tmonVFeHmVos2edlKix0X5Mjkbw9qHN4KCyCXlC
7xDB0uRX7XJIU3BGQPtUX8qEmRLE9LdizNYiRYuQfBMsUHGPgVMzppZj651G7vghOrO6E0Ga9k/U
/4sFZs0IORmtqB3EFAUO3TBXn6WN7+BfFwk3DlTNsitnpsR2iqQlb/TBwt1a/6F1cDpYB+z23yX1
27iCmYTyCebDKZQ3YytokBRW9RPlEY7v+VHuR+aL64/p7kbcJRE51CpajBJMRxU9RLGc6aF1966g
fm+QxpJJokpUfE5iQTIqafenXJmvbKAxCVg4HB/3tmm4tAhrcnnohyJcy12FyPnlnH6UIVYiqc7q
JQkk1xfOYAd4sk/7F0uQzDvryRwdIsWCl2H86dZPOkCB1C1ciLGyBwpZDUCaivIq6ZdzwoQ+7JUJ
O4t9998wZ6617BbWRLyV/f1qSMqJHRxgYposEBKJCsDEeyU+bTmOMO35V+jxrVwNTGp7pgnSOSDb
xqP/IbUh+yEjV2kvOduMPUYc32Pa7O7Yno84tHqk/wd5wxaQRqaBDrfwydWut8/l96S2nzTLbJie
FmpFYmaHNuwtZdGEyWRSvzDEYygUncinPp6drwjiXe7PAajz7vML4lpy3kMRAffEniF/nEU7A06n
UN1PAylKhcvYEiiMX5qJkGmDXWYboq7yKj+G7HsAzDoOnKCLVwTIRzAY+oRe2IlMGeOdLYt6wpgd
VtdnUaNozcd8oUAvRZuC1wfhrZQc1JgByQQnsanK7flSgdIs6PG/UySPyh3tsQVAmSSQ5HN9Bkdt
+yDnp7Ri8Q0rj/aAqBzVBJ9IVz488rk01h8P9e3XvVbGBUxbpW5HVywO24NxQTotCpz/5K1LdXwr
o9IJoQT56i+QA2+PScLJnq3FMQKK/9kff6/EcR/pUkVV1flqyfjjYh+39z4HIQ2qpmCbG933Ohq6
CPWYFV3vyugDlcnbE3Tclh7mtZD/UCnEdoaPzwp/6Dr0oeaEbuGHZ+OItgHRdS4zD3rvU8ntE8qc
R82U3OFLCaWZdCyrLv4ZUVZFE2a5ETC9aDcPaaw39F5t/J8pZ3FVXLP6NeSb8DwdAtG4/QVrOFkn
FYXaFz+osev032c4nQlUDqPuqOVPWXoFXSP0tr+Hhksv9ETfWbpEphh3YRgJXPS7vpUKGk9UzyD8
gHe6I9xt1DenXanTSDiNC2MsrZ0NoFOV4XtDSpc2F5eh87tMlUTtDOPzuhtSuT4y6ydTUZN6Hd5e
zjTuNBY25pb743wNWoKqYMMYTITGjwbygbvCCvJE1IrQtoH7KSGQXkZJUHG+ndE82RQsj14tlMql
IfACLlp1MqAW48nT/Lb4tYDeDg0qSuk5qTSxHrEvapHTaUeuEBrNAZBG/zKmoPZjypJLBphnshw4
ga1Q8N5nZSBCn6BzYFTFJFtXe3vvU+teYOuiGflFnbEekkFG13FHVK/1DYTmKoYLymsTy74jsNOg
dhVmx27UBx29L6vYKNO/qEy3S1c/TkB97sCDPErwrdDj7kHU/OS1k+3Uc7EcH4h1w7ybvwBGdLlo
w8x3NXxLrbzNVkv6o+ns4Fi/+gJLfZ9UbV+kj2sZY8mnd4IDN8Zoo66G+6CCNbCMJg3RBm86Koyn
4h6AUuYe23l9EnJtHevtt+cDeup2vL61LtJsR56zy7gZZo5I+DgAJUzasksSlr2dLmsKhh/TEArz
sI3tNDNBFV9nJVBxOCxRI2+jHX4Z1CP/C2P0T3OeslLj2KpLc/ke69O5w3syrTcW2YsVKEqWdo1r
plYhyMjD0A1RPakjcOMPOAOSB9gviC5O3n7ukmGtx5riGORIN9mjcDegD4Y+R/KK+dk3KW6DotiI
Rkel/Ahmq70HKY+tu/UNqRPraUVNyY4R8kq8iEhOWDGf0UEHB7KyNmFpPHS7xDaoMBdNUSq5Vun0
VEeqBKdzScmPhP7TcdzwSH6R6wqsR/Gdof2CRG9f2Ah7N2O9rCRwF7Xulv1emH55qxjybVGT2i03
k6M8rGDtENhxu04h5PLBSVwAuL7zHH7/H1GP2nJD69R8ZLZyvYF0sxD8LXDopbqWsKbTHv5fwd0O
eEdESB9ywNcICdnE/QVW8KrFmMOv93e10pokGQiCz4xz77nbT1PVJ2eI1dWUxAuj75iW+wCUSGuF
Y89NZej2U5MnAkZPVnolAWuhsRMX1AlLz+wCBheQqq7Db2k+qH25ot5HMHYMEwW0XJmDAFV6HnN+
jySBk+OxZhZlSnns9l/uOleOvWwCopZglBzh5CzvD7Mqw5KYWQo3Wk+xnzdtqKSuECcHSpVtLvf8
TDFDSJ0A/1kDk7VeMW0Lg7EjrxXOxuCZBjWtoyYmEXLC0U3nmlprExS3E2l7IyuNSvD+XuXyxOu7
bldE53NrbCoQxUUK3ImqW+PCbMiH9AUkJRY7RW270PaHpRsBRDt8h814kJa7lWt5tvDWQ0imxDlu
Le2cBkgoPda7LsxbN7kXCl4PGB7hrga+ZRXdpOEKxpwAKm7e7IN6w0A71jxn+yKUXHQjj9GtaXuu
ehbleAryYZh969c87gwfjnm7nnFtpzT0r+6fv0eR5L1FC49WD9pXu9HBQ3nDwKd5wvq5B+1kuyLU
Be+vqTXs2VjK6PZFR5zk6jg9m8Aa+8mGtKc6PDz0qaEVygoE3jFls6GlpLEUO4GGaykXltxm4Mdo
18n+bwLq2JjHp6wL7wsykhrh/addsj/737RrtDxhnIBiqmFWYjjy2AzS0+j2/DiLndf5LHR5z9Tq
LIKp+yKGvTG3Odeg5h48LL9Edn2htbHd3vR7vr+elcVjXXbOy1jYzkKifIXFWXNI8pVk80sY6VfN
3iGGC2fRwVTeLzN/6oSZYdm2/9n9K6UJEvbrYyDRnlDiNUrode2hkHk9m/dCemo/5tHHCtdttveq
4Q0j
`protect end_protected
